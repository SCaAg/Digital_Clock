`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/09/02 19:21:55
// Design Name: 
// Module Name: oledDraw
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module oledDrawv2(
    input clk,
    input reset_n,
    input send_done,
    input is_draw,
    output reg spi_send,
    output reg [7:0] spi_data,
    output reg dc
    );
    reg[7:0] oled_show_buffer[8*128-1:0];//显存
    reg[7:0] oled_show_line_buffer[8*128-1:0];
    reg[9:0] counter;
    reg[3:0] cur_st;
    reg [3:0] draw_st;
    localparam WAITE=0,DRAW=1,FINISH=2;
    localparam DRAW_INIT1=0,DRAW_INIT2=1,DRAW_INIT3=2,DRAW_INIT_FINISHED=3;
    integer i;
    integer x=10,y=10;
    localparam DRAW_CLOCK=0,DRAW_LINE=1;
    reg[3:0] show_st;

    reg[25:0] fenpingCounter;
    localparam fenpingM=5000000;
    //localparam fenpingM=3;
    reg[31:0] number;

    wire clk1Hz;    

    always @(posedge clk)
        begin
        if(!reset_n)
            begin
                fenpingCounter<=0;
                number<=0;
            end
        if(fenpingCounter<fenpingM)
            fenpingCounter<=fenpingCounter+1;
        else 
            fenpingCounter<=0;
        if(clk1Hz)
            number<=number+1;
        end
          
    assign clk1Hz=(fenpingCounter==fenpingM)? 1'b1:1'b0;


    always@(posedge clk)begin
        if(!reset_n)begin
            cur_st<=WAITE;
            counter<=0;
            draw_st<=DRAW_INIT1;
            show_st<=DRAW_CLOCK;
            oled_show_buffer[0]<=8'B0000000000;
            oled_show_buffer[1]<=8'B0000000000;oled_show_buffer[2]<=8'B0000000000;oled_show_buffer[3]<=8'B0000000000;oled_show_buffer[4]<=8'B0000000000;oled_show_buffer[5]<=8'B0000000000;oled_show_buffer[6]<=8'B0000000000;oled_show_buffer[7]<=8'B0000000000;oled_show_buffer[8]<=8'B0000000000;oled_show_buffer[9]<=8'B0000000000;oled_show_buffer[10]<=8'B0000000000;oled_show_buffer[11]<=8'B0000000000;oled_show_buffer[12]<=8'B0000000000;oled_show_buffer[13]<=8'B0000000000;oled_show_buffer[14]<=8'B0000000000;oled_show_buffer[15]<=8'B0000000000;oled_show_buffer[16]<=8'B0000000000;oled_show_buffer[17]<=8'B0000000000;oled_show_buffer[18]<=8'B0000000000;oled_show_buffer[19]<=8'B0000000000;oled_show_buffer[20]<=8'B0000000000;oled_show_buffer[21]<=8'B0000000000;oled_show_buffer[22]<=8'B0000000000;oled_show_buffer[23]<=8'B0000000000;oled_show_buffer[24]<=8'B0000000000;oled_show_buffer[25]<=8'B0000000000;oled_show_buffer[26]<=8'B0000000000;oled_show_buffer[27]<=8'B0000000000;oled_show_buffer[28]<=8'B0000000000;oled_show_buffer[29]<=8'B0000000000;oled_show_buffer[30]<=8'B0000000000;oled_show_buffer[31]<=8'B0000000000;oled_show_buffer[32]<=8'B0000000000;oled_show_buffer[33]<=8'B0000000000;oled_show_buffer[34]<=8'B0000000000;oled_show_buffer[35]<=8'B0000000000;oled_show_buffer[36]<=8'B0000000000;oled_show_buffer[37]<=8'B0000000000;oled_show_buffer[38]<=8'B0000000000;oled_show_buffer[39]<=8'B0000000000;oled_show_buffer[40]<=8'B0000000000;oled_show_buffer[41]<=8'B0000000000;oled_show_buffer[42]<=8'B0000000000;oled_show_buffer[43]<=8'B0000000000;oled_show_buffer[44]<=8'B0000000000;oled_show_buffer[45]<=8'B0000000000;oled_show_buffer[46]<=8'B0000000000;oled_show_buffer[47]<=8'B0010000000;oled_show_buffer[48]<=8'B0001000000;oled_show_buffer[49]<=8'B0000100000;oled_show_buffer[50]<=8'B0000100000;oled_show_buffer[51]<=8'B0011010000;oled_show_buffer[52]<=8'B0000010000;oled_show_buffer[53]<=8'B0000001000;oled_show_buffer[54]<=8'B0000001000;oled_show_buffer[55]<=8'B0000001000;oled_show_buffer[56]<=8'B0000000100;oled_show_buffer[57]<=8'B0000000100;oled_show_buffer[58]<=8'B0000000100;oled_show_buffer[59]<=8'B0000000100;oled_show_buffer[60]<=8'B0000000010;oled_show_buffer[61]<=8'B0000000010;oled_show_buffer[62]<=8'B0000000010;oled_show_buffer[63]<=8'B0000000010;oled_show_buffer[64]<=8'B0000011110;oled_show_buffer[65]<=8'B0000000010;oled_show_buffer[66]<=8'B0000000010;oled_show_buffer[67]<=8'B0000000010;oled_show_buffer[68]<=8'B0000000010;oled_show_buffer[69]<=8'B0000000010;oled_show_buffer[70]<=8'B0000000100;oled_show_buffer[71]<=8'B0000000100;oled_show_buffer[72]<=8'B0000000100;oled_show_buffer[73]<=8'B0000000100;oled_show_buffer[74]<=8'B0000001000;oled_show_buffer[75]<=8'B0000001000;oled_show_buffer[76]<=8'B0000001000;oled_show_buffer[77]<=8'B0000010000;oled_show_buffer[78]<=8'B0010010000;oled_show_buffer[79]<=8'B0001100000;oled_show_buffer[80]<=8'B0000100000;oled_show_buffer[81]<=8'B0001000000;oled_show_buffer[82]<=8'B0010000000;oled_show_buffer[83]<=8'B0000000000;oled_show_buffer[84]<=8'B0000000000;oled_show_buffer[85]<=8'B0000000000;oled_show_buffer[86]<=8'B0000000000;oled_show_buffer[87]<=8'B0000000000;oled_show_buffer[88]<=8'B0000000000;oled_show_buffer[89]<=8'B0000000000;oled_show_buffer[90]<=8'B0000000000;oled_show_buffer[91]<=8'B0000000000;oled_show_buffer[92]<=8'B0000000000;oled_show_buffer[93]<=8'B0000000000;oled_show_buffer[94]<=8'B0000000000;oled_show_buffer[95]<=8'B0000000000;oled_show_buffer[96]<=8'B0000000000;oled_show_buffer[97]<=8'B0000000000;oled_show_buffer[98]<=8'B0000000000;oled_show_buffer[99]<=8'B0000000000;oled_show_buffer[100]<=8'B0000000000;oled_show_buffer[101]<=8'B0000000000;oled_show_buffer[102]<=8'B0000000000;oled_show_buffer[103]<=8'B0000000000;oled_show_buffer[104]<=8'B0000000000;oled_show_buffer[105]<=8'B0000000000;oled_show_buffer[106]<=8'B0000000000;oled_show_buffer[107]<=8'B0000000000;oled_show_buffer[108]<=8'B0000000000;oled_show_buffer[109]<=8'B0000000000;oled_show_buffer[110]<=8'B0000000000;oled_show_buffer[111]<=8'B0000000000;oled_show_buffer[112]<=8'B0000000000;oled_show_buffer[113]<=8'B0000000000;oled_show_buffer[114]<=8'B0000000000;oled_show_buffer[115]<=8'B0000000000;oled_show_buffer[116]<=8'B0000000000;oled_show_buffer[117]<=8'B0000000000;oled_show_buffer[118]<=8'B0000000000;oled_show_buffer[119]<=8'B0000000000;oled_show_buffer[120]<=8'B0000000000;oled_show_buffer[121]<=8'B0000000000;oled_show_buffer[122]<=8'B0000000000;oled_show_buffer[123]<=8'B0000000000;oled_show_buffer[124]<=8'B0000000000;oled_show_buffer[125]<=8'B0000000000;oled_show_buffer[126]<=8'B0000000000;oled_show_buffer[127]<=8'B0000000000;oled_show_buffer[128]<=8'B0000000000;
            oled_show_buffer[129]<=8'B0000000000;oled_show_buffer[130]<=8'B0000000000;oled_show_buffer[131]<=8'B0000000000;oled_show_buffer[132]<=8'B0000000000;oled_show_buffer[133]<=8'B0000000000;oled_show_buffer[134]<=8'B0000000000;oled_show_buffer[135]<=8'B0000000000;oled_show_buffer[136]<=8'B0000000000;oled_show_buffer[137]<=8'B0000000000;oled_show_buffer[138]<=8'B0000000000;oled_show_buffer[139]<=8'B0000000000;oled_show_buffer[140]<=8'B0000000000;oled_show_buffer[141]<=8'B0000000000;oled_show_buffer[142]<=8'B0000000000;oled_show_buffer[143]<=8'B0000000000;oled_show_buffer[144]<=8'B0000000000;oled_show_buffer[145]<=8'B0000000000;oled_show_buffer[146]<=8'B0000000000;oled_show_buffer[147]<=8'B0000000000;oled_show_buffer[148]<=8'B0000000000;oled_show_buffer[149]<=8'B0000000000;oled_show_buffer[150]<=8'B0000000000;oled_show_buffer[151]<=8'B0000000000;oled_show_buffer[152]<=8'B0000000000;oled_show_buffer[153]<=8'B0000000000;oled_show_buffer[154]<=8'B0000000000;oled_show_buffer[155]<=8'B0000000000;oled_show_buffer[156]<=8'B0000000000;oled_show_buffer[157]<=8'B0000000000;oled_show_buffer[158]<=8'B0000000000;oled_show_buffer[159]<=8'B0000000000;oled_show_buffer[160]<=8'B0000000000;oled_show_buffer[161]<=8'B0000000000;oled_show_buffer[162]<=8'B0000000000;oled_show_buffer[163]<=8'B0000000000;oled_show_buffer[164]<=8'B0000000000;oled_show_buffer[165]<=8'B0000000000;oled_show_buffer[166]<=8'B0000000000;oled_show_buffer[167]<=8'B0010000000;oled_show_buffer[168]<=8'B0001000000;oled_show_buffer[169]<=8'B0000110000;oled_show_buffer[170]<=8'B0000001000;oled_show_buffer[171]<=8'B0000000100;oled_show_buffer[172]<=8'B0000000010;oled_show_buffer[173]<=8'B0000000001;oled_show_buffer[174]<=8'B0000000001;oled_show_buffer[175]<=8'B0000000000;oled_show_buffer[176]<=8'B0000000000;oled_show_buffer[177]<=8'B0000000000;oled_show_buffer[178]<=8'B0000000000;oled_show_buffer[179]<=8'B0000000000;oled_show_buffer[180]<=8'B0000000011;oled_show_buffer[181]<=8'B0000000100;oled_show_buffer[182]<=8'B0000000000;oled_show_buffer[183]<=8'B0000000000;oled_show_buffer[184]<=8'B0000000000;oled_show_buffer[185]<=8'B0000000000;oled_show_buffer[186]<=8'B0000000000;oled_show_buffer[187]<=8'B0000000000;oled_show_buffer[188]<=8'B0000000000;oled_show_buffer[189]<=8'B0000000000;oled_show_buffer[190]<=8'B0000000000;oled_show_buffer[191]<=8'B0000000000;oled_show_buffer[192]<=8'B0000000000;oled_show_buffer[193]<=8'B0000000000;oled_show_buffer[194]<=8'B0000000000;oled_show_buffer[195]<=8'B0000000000;oled_show_buffer[196]<=8'B0000000000;oled_show_buffer[197]<=8'B0000000000;oled_show_buffer[198]<=8'B0000000000;oled_show_buffer[199]<=8'B0000000000;oled_show_buffer[200]<=8'B0000000000;oled_show_buffer[201]<=8'B0000000000;oled_show_buffer[202]<=8'B0000000000;oled_show_buffer[203]<=8'B0000000000;oled_show_buffer[204]<=8'B0000000100;oled_show_buffer[205]<=8'B0000000011;oled_show_buffer[206]<=8'B0000000000;oled_show_buffer[207]<=8'B0000000000;oled_show_buffer[208]<=8'B0000000000;oled_show_buffer[209]<=8'B0000000000;oled_show_buffer[210]<=8'B0000000000;oled_show_buffer[211]<=8'B0000000001;oled_show_buffer[212]<=8'B0000000001;oled_show_buffer[213]<=8'B0000000010;oled_show_buffer[214]<=8'B0000000100;oled_show_buffer[215]<=8'B0000001000;oled_show_buffer[216]<=8'B0000110000;oled_show_buffer[217]<=8'B0001000000;oled_show_buffer[218]<=8'B0010000000;oled_show_buffer[219]<=8'B0000000000;oled_show_buffer[220]<=8'B0000000000;oled_show_buffer[221]<=8'B0000000000;oled_show_buffer[222]<=8'B0000000000;oled_show_buffer[223]<=8'B0000000000;oled_show_buffer[224]<=8'B0000000000;oled_show_buffer[225]<=8'B0000000000;oled_show_buffer[226]<=8'B0000000000;oled_show_buffer[227]<=8'B0000000000;oled_show_buffer[228]<=8'B0000000000;oled_show_buffer[229]<=8'B0000000000;oled_show_buffer[230]<=8'B0000000000;oled_show_buffer[231]<=8'B0000000000;oled_show_buffer[232]<=8'B0000000000;oled_show_buffer[233]<=8'B0000000000;oled_show_buffer[234]<=8'B0000000000;oled_show_buffer[235]<=8'B0000000000;oled_show_buffer[236]<=8'B0000000000;oled_show_buffer[237]<=8'B0000000000;oled_show_buffer[238]<=8'B0000000000;oled_show_buffer[239]<=8'B0000000000;oled_show_buffer[240]<=8'B0000000000;oled_show_buffer[241]<=8'B0000000000;oled_show_buffer[242]<=8'B0000000000;oled_show_buffer[243]<=8'B0000000000;oled_show_buffer[244]<=8'B0000000000;oled_show_buffer[245]<=8'B0000000000;oled_show_buffer[246]<=8'B0000000000;oled_show_buffer[247]<=8'B0000000000;oled_show_buffer[248]<=8'B0000000000;oled_show_buffer[249]<=8'B0000000000;oled_show_buffer[250]<=8'B0000000000;oled_show_buffer[251]<=8'B0000000000;oled_show_buffer[252]<=8'B0000000000;oled_show_buffer[253]<=8'B0000000000;oled_show_buffer[254]<=8'B0000000000;oled_show_buffer[255]<=8'B0000000000;oled_show_buffer[256]<=8'B0000000000;
            oled_show_buffer[257]<=8'B0000000000;oled_show_buffer[258]<=8'B0000000000;oled_show_buffer[259]<=8'B0000000000;oled_show_buffer[260]<=8'B0000000000;oled_show_buffer[261]<=8'B0000000000;oled_show_buffer[262]<=8'B0000000000;oled_show_buffer[263]<=8'B0000000000;oled_show_buffer[264]<=8'B0000000000;oled_show_buffer[265]<=8'B0000000000;oled_show_buffer[266]<=8'B0000000000;oled_show_buffer[267]<=8'B0000000000;oled_show_buffer[268]<=8'B0000000000;oled_show_buffer[269]<=8'B0000000000;oled_show_buffer[270]<=8'B0000000000;oled_show_buffer[271]<=8'B0000000000;oled_show_buffer[272]<=8'B0000000000;oled_show_buffer[273]<=8'B0000000000;oled_show_buffer[274]<=8'B0000000000;oled_show_buffer[275]<=8'B0000000000;oled_show_buffer[276]<=8'B0000000000;oled_show_buffer[277]<=8'B0000000000;oled_show_buffer[278]<=8'B0000000000;oled_show_buffer[279]<=8'B0000000000;oled_show_buffer[280]<=8'B0000000000;oled_show_buffer[281]<=8'B0000000000;oled_show_buffer[282]<=8'B0000000000;oled_show_buffer[283]<=8'B0000000000;oled_show_buffer[284]<=8'B0000000000;oled_show_buffer[285]<=8'B0000000000;oled_show_buffer[286]<=8'B0000000000;oled_show_buffer[287]<=8'B0000000000;oled_show_buffer[288]<=8'B0000000000;oled_show_buffer[289]<=8'B0000000000;oled_show_buffer[290]<=8'B0000000000;oled_show_buffer[291]<=8'B0010000000;oled_show_buffer[292]<=8'B0001110000;oled_show_buffer[293]<=8'B0000001100;oled_show_buffer[294]<=8'B0000000011;oled_show_buffer[295]<=8'B0000000100;oled_show_buffer[296]<=8'B0000000100;oled_show_buffer[297]<=8'B0000001000;oled_show_buffer[298]<=8'B0000001000;oled_show_buffer[299]<=8'B0000010000;oled_show_buffer[300]<=8'B0000000000;oled_show_buffer[301]<=8'B0000000000;oled_show_buffer[302]<=8'B0000000000;oled_show_buffer[303]<=8'B0000000000;oled_show_buffer[304]<=8'B0000000000;oled_show_buffer[305]<=8'B0000000000;oled_show_buffer[306]<=8'B0000000000;oled_show_buffer[307]<=8'B0000000000;oled_show_buffer[308]<=8'B0000000000;oled_show_buffer[309]<=8'B0000000000;oled_show_buffer[310]<=8'B0000000000;oled_show_buffer[311]<=8'B0000000000;oled_show_buffer[312]<=8'B0000000000;oled_show_buffer[313]<=8'B0000000000;oled_show_buffer[314]<=8'B0000000000;oled_show_buffer[315]<=8'B0000000000;oled_show_buffer[316]<=8'B0000000000;oled_show_buffer[317]<=8'B0000000000;oled_show_buffer[318]<=8'B0000000000;oled_show_buffer[319]<=8'B0000000000;oled_show_buffer[320]<=8'B0000000000;oled_show_buffer[321]<=8'B0000000000;oled_show_buffer[322]<=8'B0000000000;oled_show_buffer[323]<=8'B0000000000;oled_show_buffer[324]<=8'B0000000000;oled_show_buffer[325]<=8'B0000000000;oled_show_buffer[326]<=8'B0000000000;oled_show_buffer[327]<=8'B0000000000;oled_show_buffer[328]<=8'B0000000000;oled_show_buffer[329]<=8'B0000000000;oled_show_buffer[330]<=8'B0000000000;oled_show_buffer[331]<=8'B0000000000;oled_show_buffer[332]<=8'B0000000000;oled_show_buffer[333]<=8'B0000000000;oled_show_buffer[334]<=8'B0000000000;oled_show_buffer[335]<=8'B0000000000;oled_show_buffer[336]<=8'B0000000000;oled_show_buffer[337]<=8'B0000000000;oled_show_buffer[338]<=8'B0000000000;oled_show_buffer[339]<=8'B0000000000;oled_show_buffer[340]<=8'B0000000000;oled_show_buffer[341]<=8'B0000000000;oled_show_buffer[342]<=8'B0000100000;oled_show_buffer[343]<=8'B0000010000;oled_show_buffer[344]<=8'B0000010000;oled_show_buffer[345]<=8'B0000001000;oled_show_buffer[346]<=8'B0000001000;oled_show_buffer[347]<=8'B0000000111;oled_show_buffer[348]<=8'B0000001100;oled_show_buffer[349]<=8'B0001110000;oled_show_buffer[350]<=8'B0010000000;oled_show_buffer[351]<=8'B0000000000;oled_show_buffer[352]<=8'B0000000000;oled_show_buffer[353]<=8'B0000000000;oled_show_buffer[354]<=8'B0000000000;oled_show_buffer[355]<=8'B0000000000;oled_show_buffer[356]<=8'B0000000000;oled_show_buffer[357]<=8'B0000000000;oled_show_buffer[358]<=8'B0000000000;oled_show_buffer[359]<=8'B0000000000;oled_show_buffer[360]<=8'B0000000000;oled_show_buffer[361]<=8'B0000000000;oled_show_buffer[362]<=8'B0000000000;oled_show_buffer[363]<=8'B0000000000;oled_show_buffer[364]<=8'B0000000000;oled_show_buffer[365]<=8'B0000000000;oled_show_buffer[366]<=8'B0000000000;oled_show_buffer[367]<=8'B0000000000;oled_show_buffer[368]<=8'B0000000000;oled_show_buffer[369]<=8'B0000000000;oled_show_buffer[370]<=8'B0000000000;oled_show_buffer[371]<=8'B0000000000;oled_show_buffer[372]<=8'B0000000000;oled_show_buffer[373]<=8'B0000000000;oled_show_buffer[374]<=8'B0000000000;oled_show_buffer[375]<=8'B0000000000;oled_show_buffer[376]<=8'B0000000000;oled_show_buffer[377]<=8'B0000000000;oled_show_buffer[378]<=8'B0000000000;oled_show_buffer[379]<=8'B0000000000;oled_show_buffer[380]<=8'B0000000000;oled_show_buffer[381]<=8'B0000000000;oled_show_buffer[382]<=8'B0000000000;oled_show_buffer[383]<=8'B0000000000;oled_show_buffer[384]<=8'B0000000000;
            oled_show_buffer[385]<=8'B0000000000;oled_show_buffer[386]<=8'B0000000000;oled_show_buffer[387]<=8'B0000000000;oled_show_buffer[388]<=8'B0000000000;oled_show_buffer[389]<=8'B0000000000;oled_show_buffer[390]<=8'B0000000000;oled_show_buffer[391]<=8'B0000000000;oled_show_buffer[392]<=8'B0000000000;oled_show_buffer[393]<=8'B0000000000;oled_show_buffer[394]<=8'B0000000000;oled_show_buffer[395]<=8'B0000000000;oled_show_buffer[396]<=8'B0000000000;oled_show_buffer[397]<=8'B0000000000;oled_show_buffer[398]<=8'B0000000000;oled_show_buffer[399]<=8'B0000000000;oled_show_buffer[400]<=8'B0000000000;oled_show_buffer[401]<=8'B0000000000;oled_show_buffer[402]<=8'B0000000000;oled_show_buffer[403]<=8'B0000000000;oled_show_buffer[404]<=8'B0000000000;oled_show_buffer[405]<=8'B0000000000;oled_show_buffer[406]<=8'B0000000000;oled_show_buffer[407]<=8'B0000000000;oled_show_buffer[408]<=8'B0000000000;oled_show_buffer[409]<=8'B0000000000;oled_show_buffer[410]<=8'B0000000000;oled_show_buffer[411]<=8'B0000000000;oled_show_buffer[412]<=8'B0000000000;oled_show_buffer[413]<=8'B0000000000;oled_show_buffer[414]<=8'B0000000000;oled_show_buffer[415]<=8'B0000000000;oled_show_buffer[416]<=8'B0000000000;oled_show_buffer[417]<=8'B0000000000;oled_show_buffer[418]<=8'B0011111000;oled_show_buffer[419]<=8'B0000000111;oled_show_buffer[420]<=8'B0000000000;oled_show_buffer[421]<=8'B0000000000;oled_show_buffer[422]<=8'B0000000000;oled_show_buffer[423]<=8'B0000000000;oled_show_buffer[424]<=8'B0000000000;oled_show_buffer[425]<=8'B0000000000;oled_show_buffer[426]<=8'B0000000000;oled_show_buffer[427]<=8'B0000000000;oled_show_buffer[428]<=8'B0000000000;oled_show_buffer[429]<=8'B0000000000;oled_show_buffer[430]<=8'B0000000000;oled_show_buffer[431]<=8'B0000000000;oled_show_buffer[432]<=8'B0000000000;oled_show_buffer[433]<=8'B0000000000;oled_show_buffer[434]<=8'B0000000000;oled_show_buffer[435]<=8'B0000000000;oled_show_buffer[436]<=8'B0000000000;oled_show_buffer[437]<=8'B0000000000;oled_show_buffer[438]<=8'B0000000000;oled_show_buffer[439]<=8'B0000000000;oled_show_buffer[440]<=8'B0000000000;oled_show_buffer[441]<=8'B0000000000;oled_show_buffer[442]<=8'B0000000000;oled_show_buffer[443]<=8'B0000000000;oled_show_buffer[444]<=8'B0000000000;oled_show_buffer[445]<=8'B0000000000;oled_show_buffer[446]<=8'B0000000000;oled_show_buffer[447]<=8'B0010000000;oled_show_buffer[448]<=8'B0010000000;oled_show_buffer[449]<=8'B0010000000;oled_show_buffer[450]<=8'B0000000000;oled_show_buffer[451]<=8'B0000000000;oled_show_buffer[452]<=8'B0000000000;oled_show_buffer[453]<=8'B0000000000;oled_show_buffer[454]<=8'B0000000000;oled_show_buffer[455]<=8'B0000000000;oled_show_buffer[456]<=8'B0000000000;oled_show_buffer[457]<=8'B0000000000;oled_show_buffer[458]<=8'B0000000000;oled_show_buffer[459]<=8'B0000000000;oled_show_buffer[460]<=8'B0000000000;oled_show_buffer[461]<=8'B0000000000;oled_show_buffer[462]<=8'B0000000000;oled_show_buffer[463]<=8'B0000000000;oled_show_buffer[464]<=8'B0000000000;oled_show_buffer[465]<=8'B0000000000;oled_show_buffer[466]<=8'B0000000000;oled_show_buffer[467]<=8'B0000000000;oled_show_buffer[468]<=8'B0000000000;oled_show_buffer[469]<=8'B0000000000;oled_show_buffer[470]<=8'B0000000000;oled_show_buffer[471]<=8'B0000000000;oled_show_buffer[472]<=8'B0000000000;oled_show_buffer[473]<=8'B0000000000;oled_show_buffer[474]<=8'B0000000000;oled_show_buffer[475]<=8'B0000000000;oled_show_buffer[476]<=8'B0000000000;oled_show_buffer[477]<=8'B0000000000;oled_show_buffer[478]<=8'B0000000111;oled_show_buffer[479]<=8'B0011111000;oled_show_buffer[480]<=8'B0000000000;oled_show_buffer[481]<=8'B0000000000;oled_show_buffer[482]<=8'B0000000000;oled_show_buffer[483]<=8'B0000000000;oled_show_buffer[484]<=8'B0000000000;oled_show_buffer[485]<=8'B0000000000;oled_show_buffer[486]<=8'B0000000000;oled_show_buffer[487]<=8'B0000000000;oled_show_buffer[488]<=8'B0000000000;oled_show_buffer[489]<=8'B0000000000;oled_show_buffer[490]<=8'B0000000000;oled_show_buffer[491]<=8'B0000000000;oled_show_buffer[492]<=8'B0000000000;oled_show_buffer[493]<=8'B0000000000;oled_show_buffer[494]<=8'B0000000000;oled_show_buffer[495]<=8'B0000000000;oled_show_buffer[496]<=8'B0000000000;oled_show_buffer[497]<=8'B0000000000;oled_show_buffer[498]<=8'B0000000000;oled_show_buffer[499]<=8'B0000000000;oled_show_buffer[500]<=8'B0000000000;oled_show_buffer[501]<=8'B0000000000;oled_show_buffer[502]<=8'B0000000000;oled_show_buffer[503]<=8'B0000000000;oled_show_buffer[504]<=8'B0000000000;oled_show_buffer[505]<=8'B0000000000;oled_show_buffer[506]<=8'B0000000000;oled_show_buffer[507]<=8'B0000000000;oled_show_buffer[508]<=8'B0000000000;oled_show_buffer[509]<=8'B0000000000;oled_show_buffer[510]<=8'B0000000000;oled_show_buffer[511]<=8'B0000000000;oled_show_buffer[512]<=8'B0000000000;
            oled_show_buffer[513]<=8'B0000000000;oled_show_buffer[514]<=8'B0000000000;oled_show_buffer[515]<=8'B0000000000;oled_show_buffer[516]<=8'B0000000000;oled_show_buffer[517]<=8'B0000000000;oled_show_buffer[518]<=8'B0000000000;oled_show_buffer[519]<=8'B0000000000;oled_show_buffer[520]<=8'B0000000000;oled_show_buffer[521]<=8'B0000000000;oled_show_buffer[522]<=8'B0000000000;oled_show_buffer[523]<=8'B0000000000;oled_show_buffer[524]<=8'B0000000000;oled_show_buffer[525]<=8'B0000000000;oled_show_buffer[526]<=8'B0000000000;oled_show_buffer[527]<=8'B0000000000;oled_show_buffer[528]<=8'B0000000000;oled_show_buffer[529]<=8'B0000000000;oled_show_buffer[530]<=8'B0000000000;oled_show_buffer[531]<=8'B0000000000;oled_show_buffer[532]<=8'B0000000010;oled_show_buffer[533]<=8'B0000000000;oled_show_buffer[534]<=8'B0000000000;oled_show_buffer[535]<=8'B0000000000;oled_show_buffer[536]<=8'B0000000000;oled_show_buffer[537]<=8'B0000000000;oled_show_buffer[538]<=8'B0000000000;oled_show_buffer[539]<=8'B0000000000;oled_show_buffer[540]<=8'B0000000000;oled_show_buffer[541]<=8'B0000000000;oled_show_buffer[542]<=8'B0000000000;oled_show_buffer[543]<=8'B0000000000;oled_show_buffer[544]<=8'B0000000000;oled_show_buffer[545]<=8'B0000000000;oled_show_buffer[546]<=8'B0000011111;oled_show_buffer[547]<=8'B0011100001;oled_show_buffer[548]<=8'B0000000001;oled_show_buffer[549]<=8'B0000000001;oled_show_buffer[550]<=8'B0000000001;oled_show_buffer[551]<=8'B0000000000;oled_show_buffer[552]<=8'B0000000000;oled_show_buffer[553]<=8'B0000000000;oled_show_buffer[554]<=8'B0000000000;oled_show_buffer[555]<=8'B0000000000;oled_show_buffer[556]<=8'B0000000000;oled_show_buffer[557]<=8'B0000000000;oled_show_buffer[558]<=8'B0000000000;oled_show_buffer[559]<=8'B0000000000;oled_show_buffer[560]<=8'B0000000000;oled_show_buffer[561]<=8'B0000000000;oled_show_buffer[562]<=8'B0000000000;oled_show_buffer[563]<=8'B0000000000;oled_show_buffer[564]<=8'B0000000000;oled_show_buffer[565]<=8'B0000000000;oled_show_buffer[566]<=8'B0000000000;oled_show_buffer[567]<=8'B0000000000;oled_show_buffer[568]<=8'B0000000000;oled_show_buffer[569]<=8'B0000000000;oled_show_buffer[570]<=8'B0000000000;oled_show_buffer[571]<=8'B0000000000;oled_show_buffer[572]<=8'B0000000000;oled_show_buffer[573]<=8'B0000000000;oled_show_buffer[574]<=8'B0000000000;oled_show_buffer[575]<=8'B0000000011;oled_show_buffer[576]<=8'B0000000011;oled_show_buffer[577]<=8'B0000000011;oled_show_buffer[578]<=8'B0000000000;oled_show_buffer[579]<=8'B0000000000;oled_show_buffer[580]<=8'B0000000000;oled_show_buffer[581]<=8'B0000000000;oled_show_buffer[582]<=8'B0000000000;oled_show_buffer[583]<=8'B0000000000;oled_show_buffer[584]<=8'B0000000000;oled_show_buffer[585]<=8'B0000000000;oled_show_buffer[586]<=8'B0000000000;oled_show_buffer[587]<=8'B0000000000;oled_show_buffer[588]<=8'B0000000000;oled_show_buffer[589]<=8'B0000000000;oled_show_buffer[590]<=8'B0000000000;oled_show_buffer[591]<=8'B0000000000;oled_show_buffer[592]<=8'B0000000000;oled_show_buffer[593]<=8'B0000000000;oled_show_buffer[594]<=8'B0000000000;oled_show_buffer[595]<=8'B0000000000;oled_show_buffer[596]<=8'B0000000000;oled_show_buffer[597]<=8'B0000000000;oled_show_buffer[598]<=8'B0000000000;oled_show_buffer[599]<=8'B0000000000;oled_show_buffer[600]<=8'B0000000000;oled_show_buffer[601]<=8'B0000000000;oled_show_buffer[602]<=8'B0000000000;oled_show_buffer[603]<=8'B0000000000;oled_show_buffer[604]<=8'B0000000001;oled_show_buffer[605]<=8'B0000000001;oled_show_buffer[606]<=8'B0011100001;oled_show_buffer[607]<=8'B0000011111;oled_show_buffer[608]<=8'B0000000000;oled_show_buffer[609]<=8'B0000000000;oled_show_buffer[610]<=8'B0000000000;oled_show_buffer[611]<=8'B0000000000;oled_show_buffer[612]<=8'B0000000000;oled_show_buffer[613]<=8'B0000000000;oled_show_buffer[614]<=8'B0000000000;oled_show_buffer[615]<=8'B0000000000;oled_show_buffer[616]<=8'B0000000000;oled_show_buffer[617]<=8'B0000000000;oled_show_buffer[618]<=8'B0000000000;oled_show_buffer[619]<=8'B0000000000;oled_show_buffer[620]<=8'B0000000000;oled_show_buffer[621]<=8'B0000000000;oled_show_buffer[622]<=8'B0000000000;oled_show_buffer[623]<=8'B0000000000;oled_show_buffer[624]<=8'B0000000000;oled_show_buffer[625]<=8'B0000000000;oled_show_buffer[626]<=8'B0000000000;oled_show_buffer[627]<=8'B0000000000;oled_show_buffer[628]<=8'B0000000000;oled_show_buffer[629]<=8'B0000000000;oled_show_buffer[630]<=8'B0000000000;oled_show_buffer[631]<=8'B0000000000;oled_show_buffer[632]<=8'B0000000000;oled_show_buffer[633]<=8'B0000000000;oled_show_buffer[634]<=8'B0000000000;oled_show_buffer[635]<=8'B0000000000;oled_show_buffer[636]<=8'B0000000000;oled_show_buffer[637]<=8'B0000000000;oled_show_buffer[638]<=8'B0000000000;oled_show_buffer[639]<=8'B0000000000;oled_show_buffer[640]<=8'B0000000000;
            oled_show_buffer[641]<=8'B0000000000;oled_show_buffer[642]<=8'B0000000000;oled_show_buffer[643]<=8'B0000000000;oled_show_buffer[644]<=8'B0000000000;oled_show_buffer[645]<=8'B0000000000;oled_show_buffer[646]<=8'B0000000000;oled_show_buffer[647]<=8'B0000000000;oled_show_buffer[648]<=8'B0000000000;oled_show_buffer[649]<=8'B0000000000;oled_show_buffer[650]<=8'B0000000000;oled_show_buffer[651]<=8'B0000000000;oled_show_buffer[652]<=8'B0000000000;oled_show_buffer[653]<=8'B0000000000;oled_show_buffer[654]<=8'B0000000000;oled_show_buffer[655]<=8'B0000000000;oled_show_buffer[656]<=8'B0000000000;oled_show_buffer[657]<=8'B0000000000;oled_show_buffer[658]<=8'B0000000000;oled_show_buffer[659]<=8'B0000000000;oled_show_buffer[660]<=8'B0000000000;oled_show_buffer[661]<=8'B0000000000;oled_show_buffer[662]<=8'B0000000000;oled_show_buffer[663]<=8'B0000000000;oled_show_buffer[664]<=8'B0000000000;oled_show_buffer[665]<=8'B0000000000;oled_show_buffer[666]<=8'B0000000000;oled_show_buffer[667]<=8'B0000000000;oled_show_buffer[668]<=8'B0000000000;oled_show_buffer[669]<=8'B0000000000;oled_show_buffer[670]<=8'B0000000000;oled_show_buffer[671]<=8'B0000000000;oled_show_buffer[672]<=8'B0000000000;oled_show_buffer[673]<=8'B0000000000;oled_show_buffer[674]<=8'B0000000000;oled_show_buffer[675]<=8'B0000000001;oled_show_buffer[676]<=8'B0000001110;oled_show_buffer[677]<=8'B0000110000;oled_show_buffer[678]<=8'B0011000000;oled_show_buffer[679]<=8'B0000100000;oled_show_buffer[680]<=8'B0000100000;oled_show_buffer[681]<=8'B0000010000;oled_show_buffer[682]<=8'B0000010000;oled_show_buffer[683]<=8'B0000001000;oled_show_buffer[684]<=8'B0000000000;oled_show_buffer[685]<=8'B0000000000;oled_show_buffer[686]<=8'B0000000000;oled_show_buffer[687]<=8'B0000000000;oled_show_buffer[688]<=8'B0000000000;oled_show_buffer[689]<=8'B0000000000;oled_show_buffer[690]<=8'B0000000000;oled_show_buffer[691]<=8'B0000000000;oled_show_buffer[692]<=8'B0000000000;oled_show_buffer[693]<=8'B0000000000;oled_show_buffer[694]<=8'B0000000000;oled_show_buffer[695]<=8'B0000000000;oled_show_buffer[696]<=8'B0000000000;oled_show_buffer[697]<=8'B0000000000;oled_show_buffer[698]<=8'B0000000000;oled_show_buffer[699]<=8'B0000000000;oled_show_buffer[700]<=8'B0000000000;oled_show_buffer[701]<=8'B0000000000;oled_show_buffer[702]<=8'B0000000000;oled_show_buffer[703]<=8'B0000000000;oled_show_buffer[704]<=8'B0000000000;oled_show_buffer[705]<=8'B0000000000;oled_show_buffer[706]<=8'B0000000000;oled_show_buffer[707]<=8'B0000000000;oled_show_buffer[708]<=8'B0000000000;oled_show_buffer[709]<=8'B0000000000;oled_show_buffer[710]<=8'B0000000000;oled_show_buffer[711]<=8'B0000000000;oled_show_buffer[712]<=8'B0000000000;oled_show_buffer[713]<=8'B0000000000;oled_show_buffer[714]<=8'B0000000000;oled_show_buffer[715]<=8'B0000000000;oled_show_buffer[716]<=8'B0000000000;oled_show_buffer[717]<=8'B0000000000;oled_show_buffer[718]<=8'B0000000000;oled_show_buffer[719]<=8'B0000000000;oled_show_buffer[720]<=8'B0000000000;oled_show_buffer[721]<=8'B0000000000;oled_show_buffer[722]<=8'B0000000000;oled_show_buffer[723]<=8'B0000000000;oled_show_buffer[724]<=8'B0000000000;oled_show_buffer[725]<=8'B0000001000;oled_show_buffer[726]<=8'B0000010000;oled_show_buffer[727]<=8'B0000010000;oled_show_buffer[728]<=8'B0000100000;oled_show_buffer[729]<=8'B0001000000;oled_show_buffer[730]<=8'B0001000000;oled_show_buffer[731]<=8'B0011000000;oled_show_buffer[732]<=8'B0000110000;oled_show_buffer[733]<=8'B0000001110;oled_show_buffer[734]<=8'B0000000001;oled_show_buffer[735]<=8'B0000000000;oled_show_buffer[736]<=8'B0000000000;oled_show_buffer[737]<=8'B0000000000;oled_show_buffer[738]<=8'B0000000000;oled_show_buffer[739]<=8'B0000000000;oled_show_buffer[740]<=8'B0000000000;oled_show_buffer[741]<=8'B0000000000;oled_show_buffer[742]<=8'B0000000000;oled_show_buffer[743]<=8'B0000000000;oled_show_buffer[744]<=8'B0000000000;oled_show_buffer[745]<=8'B0000000000;oled_show_buffer[746]<=8'B0000000000;oled_show_buffer[747]<=8'B0000000000;oled_show_buffer[748]<=8'B0000000000;oled_show_buffer[749]<=8'B0000000000;oled_show_buffer[750]<=8'B0000000000;oled_show_buffer[751]<=8'B0000000000;oled_show_buffer[752]<=8'B0000000000;oled_show_buffer[753]<=8'B0000000000;oled_show_buffer[754]<=8'B0000000000;oled_show_buffer[755]<=8'B0000000000;oled_show_buffer[756]<=8'B0000000000;oled_show_buffer[757]<=8'B0000000000;oled_show_buffer[758]<=8'B0000000000;oled_show_buffer[759]<=8'B0000000000;oled_show_buffer[760]<=8'B0000000000;oled_show_buffer[761]<=8'B0000000000;oled_show_buffer[762]<=8'B0000000000;oled_show_buffer[763]<=8'B0000000000;oled_show_buffer[764]<=8'B0000000000;oled_show_buffer[765]<=8'B0000000000;oled_show_buffer[766]<=8'B0000000000;oled_show_buffer[767]<=8'B0000000000;oled_show_buffer[768]<=8'B0000000000;
            oled_show_buffer[769]<=8'B0000000000;oled_show_buffer[770]<=8'B0000000000;oled_show_buffer[771]<=8'B0000000000;oled_show_buffer[772]<=8'B0000000000;oled_show_buffer[773]<=8'B0000000000;oled_show_buffer[774]<=8'B0000000000;oled_show_buffer[775]<=8'B0000000000;oled_show_buffer[776]<=8'B0000000000;oled_show_buffer[777]<=8'B0000000000;oled_show_buffer[778]<=8'B0000000000;oled_show_buffer[779]<=8'B0000000000;oled_show_buffer[780]<=8'B0000000000;oled_show_buffer[781]<=8'B0000000000;oled_show_buffer[782]<=8'B0000000000;oled_show_buffer[783]<=8'B0000000000;oled_show_buffer[784]<=8'B0000000000;oled_show_buffer[785]<=8'B0000000000;oled_show_buffer[786]<=8'B0000000000;oled_show_buffer[787]<=8'B0000000000;oled_show_buffer[788]<=8'B0000000000;oled_show_buffer[789]<=8'B0000000000;oled_show_buffer[790]<=8'B0000000000;oled_show_buffer[791]<=8'B0000000000;oled_show_buffer[792]<=8'B0000000000;oled_show_buffer[793]<=8'B0000000000;oled_show_buffer[794]<=8'B0000000000;oled_show_buffer[795]<=8'B0000000000;oled_show_buffer[796]<=8'B0000000000;oled_show_buffer[797]<=8'B0000000000;oled_show_buffer[798]<=8'B0000000000;oled_show_buffer[799]<=8'B0000000000;oled_show_buffer[800]<=8'B0000000000;oled_show_buffer[801]<=8'B0000000000;oled_show_buffer[802]<=8'B0000000000;oled_show_buffer[803]<=8'B0000000000;oled_show_buffer[804]<=8'B0000000000;oled_show_buffer[805]<=8'B0000000000;oled_show_buffer[806]<=8'B0000000000;oled_show_buffer[807]<=8'B0000000001;oled_show_buffer[808]<=8'B0000000010;oled_show_buffer[809]<=8'B0000001100;oled_show_buffer[810]<=8'B0000010000;oled_show_buffer[811]<=8'B0000100000;oled_show_buffer[812]<=8'B0001000000;oled_show_buffer[813]<=8'B0010000000;oled_show_buffer[814]<=8'B0010000000;oled_show_buffer[815]<=8'B0000000000;oled_show_buffer[816]<=8'B0000000000;oled_show_buffer[817]<=8'B0000000000;oled_show_buffer[818]<=8'B0010000000;oled_show_buffer[819]<=8'B0010000000;oled_show_buffer[820]<=8'B0001000000;oled_show_buffer[821]<=8'B0000100000;oled_show_buffer[822]<=8'B0000000000;oled_show_buffer[823]<=8'B0000000000;oled_show_buffer[824]<=8'B0000000000;oled_show_buffer[825]<=8'B0000000000;oled_show_buffer[826]<=8'B0000000000;oled_show_buffer[827]<=8'B0000000000;oled_show_buffer[828]<=8'B0000000000;oled_show_buffer[829]<=8'B0000000000;oled_show_buffer[830]<=8'B0000000000;oled_show_buffer[831]<=8'B0000000000;oled_show_buffer[832]<=8'B0000000000;oled_show_buffer[833]<=8'B0000000000;oled_show_buffer[834]<=8'B0000000000;oled_show_buffer[835]<=8'B0000000000;oled_show_buffer[836]<=8'B0000000000;oled_show_buffer[837]<=8'B0000000000;oled_show_buffer[838]<=8'B0000000000;oled_show_buffer[839]<=8'B0000000000;oled_show_buffer[840]<=8'B0000000000;oled_show_buffer[841]<=8'B0000000000;oled_show_buffer[842]<=8'B0000000000;oled_show_buffer[843]<=8'B0000000000;oled_show_buffer[844]<=8'B0001000000;oled_show_buffer[845]<=8'B0010000000;oled_show_buffer[846]<=8'B0000000000;oled_show_buffer[847]<=8'B0000000000;oled_show_buffer[848]<=8'B0000000000;oled_show_buffer[849]<=8'B0000000000;oled_show_buffer[850]<=8'B0000000000;oled_show_buffer[851]<=8'B0010000000;oled_show_buffer[852]<=8'B0010000000;oled_show_buffer[853]<=8'B0001000000;oled_show_buffer[854]<=8'B0000100000;oled_show_buffer[855]<=8'B0000010000;oled_show_buffer[856]<=8'B0000001100;oled_show_buffer[857]<=8'B0000000010;oled_show_buffer[858]<=8'B0000000001;oled_show_buffer[859]<=8'B0000000000;oled_show_buffer[860]<=8'B0000000000;oled_show_buffer[861]<=8'B0000000000;oled_show_buffer[862]<=8'B0000000000;oled_show_buffer[863]<=8'B0000000000;oled_show_buffer[864]<=8'B0000000000;oled_show_buffer[865]<=8'B0000000000;oled_show_buffer[866]<=8'B0000000000;oled_show_buffer[867]<=8'B0000000000;oled_show_buffer[868]<=8'B0000000000;oled_show_buffer[869]<=8'B0000000000;oled_show_buffer[870]<=8'B0000000000;oled_show_buffer[871]<=8'B0000000000;oled_show_buffer[872]<=8'B0000000000;oled_show_buffer[873]<=8'B0000000000;oled_show_buffer[874]<=8'B0000000000;oled_show_buffer[875]<=8'B0000000000;oled_show_buffer[876]<=8'B0000000000;oled_show_buffer[877]<=8'B0000000000;oled_show_buffer[878]<=8'B0000000000;oled_show_buffer[879]<=8'B0000000000;oled_show_buffer[880]<=8'B0000000000;oled_show_buffer[881]<=8'B0000000000;oled_show_buffer[882]<=8'B0000000000;oled_show_buffer[883]<=8'B0000000000;oled_show_buffer[884]<=8'B0000000000;oled_show_buffer[885]<=8'B0000000000;oled_show_buffer[886]<=8'B0000000000;oled_show_buffer[887]<=8'B0000000000;oled_show_buffer[888]<=8'B0000000000;oled_show_buffer[889]<=8'B0000000000;oled_show_buffer[890]<=8'B0000000000;oled_show_buffer[891]<=8'B0000000000;oled_show_buffer[892]<=8'B0000000000;oled_show_buffer[893]<=8'B0000000000;oled_show_buffer[894]<=8'B0000000000;oled_show_buffer[895]<=8'B0000000000;oled_show_buffer[896]<=8'B0000000000;
            oled_show_buffer[897]<=8'B0000000000;oled_show_buffer[898]<=8'B0000000000;oled_show_buffer[899]<=8'B0000000000;oled_show_buffer[900]<=8'B0000000000;oled_show_buffer[901]<=8'B0000000000;oled_show_buffer[902]<=8'B0000000000;oled_show_buffer[903]<=8'B0000000000;oled_show_buffer[904]<=8'B0000000000;oled_show_buffer[905]<=8'B0000000000;oled_show_buffer[906]<=8'B0000000000;oled_show_buffer[907]<=8'B0000000000;oled_show_buffer[908]<=8'B0000000000;oled_show_buffer[909]<=8'B0000000000;oled_show_buffer[910]<=8'B0000000000;oled_show_buffer[911]<=8'B0000000000;oled_show_buffer[912]<=8'B0000000000;oled_show_buffer[913]<=8'B0000000000;oled_show_buffer[914]<=8'B0000000000;oled_show_buffer[915]<=8'B0000000000;oled_show_buffer[916]<=8'B0000000000;oled_show_buffer[917]<=8'B0000000000;oled_show_buffer[918]<=8'B0000000000;oled_show_buffer[919]<=8'B0000000000;oled_show_buffer[920]<=8'B0000000000;oled_show_buffer[921]<=8'B0000000000;oled_show_buffer[922]<=8'B0000000000;oled_show_buffer[923]<=8'B0000000000;oled_show_buffer[924]<=8'B0000000000;oled_show_buffer[925]<=8'B0000000000;oled_show_buffer[926]<=8'B0000000000;oled_show_buffer[927]<=8'B0000000000;oled_show_buffer[928]<=8'B0000000000;oled_show_buffer[929]<=8'B0000000000;oled_show_buffer[930]<=8'B0000000000;oled_show_buffer[931]<=8'B0000000000;oled_show_buffer[932]<=8'B0000000000;oled_show_buffer[933]<=8'B0000000000;oled_show_buffer[934]<=8'B0000000000;oled_show_buffer[935]<=8'B0000000000;oled_show_buffer[936]<=8'B0000000000;oled_show_buffer[937]<=8'B0000000000;oled_show_buffer[938]<=8'B0000000000;oled_show_buffer[939]<=8'B0000000000;oled_show_buffer[940]<=8'B0000000000;oled_show_buffer[941]<=8'B0000000000;oled_show_buffer[942]<=8'B0000000000;oled_show_buffer[943]<=8'B0000000001;oled_show_buffer[944]<=8'B0000000010;oled_show_buffer[945]<=8'B0000000101;oled_show_buffer[946]<=8'B0000000100;oled_show_buffer[947]<=8'B0000001000;oled_show_buffer[948]<=8'B0000001000;oled_show_buffer[949]<=8'B0000010000;oled_show_buffer[950]<=8'B0000010000;oled_show_buffer[951]<=8'B0000010000;oled_show_buffer[952]<=8'B0000100000;oled_show_buffer[953]<=8'B0000100000;oled_show_buffer[954]<=8'B0000100000;oled_show_buffer[955]<=8'B0000100000;oled_show_buffer[956]<=8'B0001000000;oled_show_buffer[957]<=8'B0001000000;oled_show_buffer[958]<=8'B0001000000;oled_show_buffer[959]<=8'B0001000000;oled_show_buffer[960]<=8'B0001000000;oled_show_buffer[961]<=8'B0001111000;oled_show_buffer[962]<=8'B0001000000;oled_show_buffer[963]<=8'B0001000000;oled_show_buffer[964]<=8'B0001000000;oled_show_buffer[965]<=8'B0001000000;oled_show_buffer[966]<=8'B0000100000;oled_show_buffer[967]<=8'B0000100000;oled_show_buffer[968]<=8'B0000100000;oled_show_buffer[969]<=8'B0000100000;oled_show_buffer[970]<=8'B0000010000;oled_show_buffer[971]<=8'B0000010000;oled_show_buffer[972]<=8'B0000010000;oled_show_buffer[973]<=8'B0000001000;oled_show_buffer[974]<=8'B0000001001;oled_show_buffer[975]<=8'B0000000110;oled_show_buffer[976]<=8'B0000000100;oled_show_buffer[977]<=8'B0000000010;oled_show_buffer[978]<=8'B0000000001;oled_show_buffer[979]<=8'B0000000000;oled_show_buffer[980]<=8'B0000000000;oled_show_buffer[981]<=8'B0000000000;oled_show_buffer[982]<=8'B0000000000;oled_show_buffer[983]<=8'B0000000000;oled_show_buffer[984]<=8'B0000000000;oled_show_buffer[985]<=8'B0000000000;oled_show_buffer[986]<=8'B0000000000;oled_show_buffer[987]<=8'B0000000000;oled_show_buffer[988]<=8'B0000000000;oled_show_buffer[989]<=8'B0000000000;oled_show_buffer[990]<=8'B0000000000;oled_show_buffer[991]<=8'B0000000000;oled_show_buffer[992]<=8'B0000000000;oled_show_buffer[993]<=8'B0000000000;oled_show_buffer[994]<=8'B0000000000;oled_show_buffer[995]<=8'B0000000000;oled_show_buffer[996]<=8'B0000000000;oled_show_buffer[997]<=8'B0000000000;oled_show_buffer[998]<=8'B0000000000;oled_show_buffer[999]<=8'B0000000000;oled_show_buffer[1000]<=8'B0000000000;oled_show_buffer[1001]<=8'B0000000000;oled_show_buffer[1002]<=8'B0000000000;oled_show_buffer[1003]<=8'B0000000000;oled_show_buffer[1004]<=8'B0000000000;oled_show_buffer[1005]<=8'B0000000000;oled_show_buffer[1006]<=8'B0000000000;oled_show_buffer[1007]<=8'B0000000000;oled_show_buffer[1008]<=8'B0000000000;oled_show_buffer[1009]<=8'B0000000000;oled_show_buffer[1010]<=8'B0000000000;oled_show_buffer[1011]<=8'B0000000000;oled_show_buffer[1012]<=8'B0000000000;oled_show_buffer[1013]<=8'B0000000000;oled_show_buffer[1014]<=8'B0000000000;oled_show_buffer[1015]<=8'B0000000000;oled_show_buffer[1016]<=8'B0000000000;oled_show_buffer[1017]<=8'B0000000000;oled_show_buffer[1018]<=8'B0000000000;oled_show_buffer[1019]<=8'B0000000000;oled_show_buffer[1020]<=8'B0000000000;oled_show_buffer[1021]<=8'B0000000000;oled_show_buffer[1022]<=8'B0000000000;oled_show_buffer[1023]<=8'B0000000000; 
        end
        case(cur_st)
            WAITE:
                if(is_draw)begin
                    cur_st<=DRAW; 
                    counter<=0;
                    draw_st<=DRAW_INIT1;
                    case(show_st)
                        DRAW_CLOCK:begin
                            for(i=0;i<1024;i=i+1)begin
                                oled_show_line_buffer[i]<=0;
                            end
                        end
                        DRAW_LINE:begin
                            case(number%60)
                            0:begin oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[448]<=8'B11111111;oled_show_line_buffer[320]<=8'B11111111;oled_show_line_buffer[192]<=8'B11111111;oled_show_line_buffer[64]<=8'B10011110;end
                            1:begin oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[448]<=8'B11111111;oled_show_line_buffer[320]<=8'B10000000;oled_show_line_buffer[321]<=8'B11111111;oled_show_line_buffer[193]<=8'B11000000;oled_show_line_buffer[194]<=8'B01111111;oled_show_line_buffer[66]<=8'B11110010;end
                            2:begin oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[448]<=8'B11110000;oled_show_line_buffer[449]<=8'B10011111;oled_show_line_buffer[450]<=8'B00000001;oled_show_line_buffer[322]<=8'B11111000;oled_show_line_buffer[323]<=8'B00001111;oled_show_line_buffer[195]<=8'B11000000;oled_show_line_buffer[196]<=8'B01111110;oled_show_line_buffer[197]<=8'B00000011;oled_show_line_buffer[69]<=8'B11100010;end
                            3:begin oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[448]<=8'B11000000;oled_show_line_buffer[449]<=8'B11111000;oled_show_line_buffer[450]<=8'B00001111;oled_show_line_buffer[451]<=8'B00000001;oled_show_line_buffer[323]<=8'B11100000;oled_show_line_buffer[324]<=8'B00111100;oled_show_line_buffer[325]<=8'B00000111;oled_show_line_buffer[197]<=8'B10000000;oled_show_line_buffer[198]<=8'B11111000;oled_show_line_buffer[199]<=8'B00001111;end
                            4:begin oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[449]<=8'B11100000;oled_show_line_buffer[450]<=8'B00111100;oled_show_line_buffer[451]<=8'B00000111;oled_show_line_buffer[452]<=8'B00000001;oled_show_line_buffer[324]<=8'B11000000;oled_show_line_buffer[325]<=8'B01110000;oled_show_line_buffer[326]<=8'B00011110;oled_show_line_buffer[327]<=8'B00000011;oled_show_line_buffer[199]<=8'B10000000;oled_show_line_buffer[200]<=8'B11100000;oled_show_line_buffer[201]<=8'B00111000;oled_show_line_buffer[202]<=8'B00001111;end
                            5:begin oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[449]<=8'B11000000;oled_show_line_buffer[450]<=8'B01110000;oled_show_line_buffer[451]<=8'B00011100;oled_show_line_buffer[452]<=8'B00000111;oled_show_line_buffer[453]<=8'B00000001;oled_show_line_buffer[325]<=8'B10000000;oled_show_line_buffer[326]<=8'B11100000;oled_show_line_buffer[327]<=8'B00111000;oled_show_line_buffer[328]<=8'B00001110;oled_show_line_buffer[329]<=8'B00000011;oled_show_line_buffer[330]<=8'B00000001;oled_show_line_buffer[202]<=8'B11000000;oled_show_line_buffer[203]<=8'B01110000;oled_show_line_buffer[204]<=8'B00011100;end
                            6:begin oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[449]<=8'B11000000;oled_show_line_buffer[450]<=8'B01100000;oled_show_line_buffer[451]<=8'B00111000;oled_show_line_buffer[452]<=8'B00001100;oled_show_line_buffer[453]<=8'B00000110;oled_show_line_buffer[454]<=8'B00000011;oled_show_line_buffer[326]<=8'B10000000;oled_show_line_buffer[327]<=8'B11000000;oled_show_line_buffer[328]<=8'B01100000;oled_show_line_buffer[329]<=8'B00111000;oled_show_line_buffer[330]<=8'B00001100;oled_show_line_buffer[331]<=8'B00000111;oled_show_line_buffer[332]<=8'B00000001;oled_show_line_buffer[204]<=8'B10000100;oled_show_line_buffer[205]<=8'B11000011;oled_show_line_buffer[206]<=8'B01110000;end
                            7:begin oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[449]<=8'B10000000;oled_show_line_buffer[450]<=8'B11000000;oled_show_line_buffer[451]<=8'B01100000;oled_show_line_buffer[452]<=8'B00111000;oled_show_line_buffer[453]<=8'B00001100;oled_show_line_buffer[454]<=8'B00000110;oled_show_line_buffer[455]<=8'B00000011;oled_show_line_buffer[456]<=8'B00000001;oled_show_line_buffer[328]<=8'B10000000;oled_show_line_buffer[329]<=8'B11000000;oled_show_line_buffer[330]<=8'B01100000;oled_show_line_buffer[331]<=8'B00110000;oled_show_line_buffer[332]<=8'B00011000;oled_show_line_buffer[333]<=8'B00001110;oled_show_line_buffer[334]<=8'B00000011;oled_show_line_buffer[335]<=8'B00000001;oled_show_line_buffer[207]<=8'B10000000;oled_show_line_buffer[208]<=8'B11000000;oled_show_line_buffer[209]<=8'B01100000;end
                            8:begin oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[449]<=8'B10000000;oled_show_line_buffer[450]<=8'B11000000;oled_show_line_buffer[451]<=8'B01100000;oled_show_line_buffer[452]<=8'B00110000;oled_show_line_buffer[453]<=8'B00010000;oled_show_line_buffer[454]<=8'B00011000;oled_show_line_buffer[455]<=8'B00001100;oled_show_line_buffer[456]<=8'B00000110;oled_show_line_buffer[457]<=8'B00000011;oled_show_line_buffer[458]<=8'B00000001;oled_show_line_buffer[330]<=8'B10000000;oled_show_line_buffer[331]<=8'B11000000;oled_show_line_buffer[332]<=8'B01100000;oled_show_line_buffer[333]<=8'B00110000;oled_show_line_buffer[334]<=8'B00011000;oled_show_line_buffer[335]<=8'B00001000;oled_show_line_buffer[336]<=8'B00001100;oled_show_line_buffer[337]<=8'B00000110;oled_show_line_buffer[338]<=8'B00000011;end
                            9:begin oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[578]<=8'B00000001;oled_show_line_buffer[450]<=8'B10000000;oled_show_line_buffer[451]<=8'B11000000;oled_show_line_buffer[452]<=8'B01100000;oled_show_line_buffer[453]<=8'B00100000;oled_show_line_buffer[454]<=8'B00110000;oled_show_line_buffer[455]<=8'B00011000;oled_show_line_buffer[456]<=8'B00001100;oled_show_line_buffer[457]<=8'B00000100;oled_show_line_buffer[458]<=8'B00000110;oled_show_line_buffer[459]<=8'B00000011;oled_show_line_buffer[460]<=8'B00000001;oled_show_line_buffer[461]<=8'B00000001;oled_show_line_buffer[333]<=8'B10000000;oled_show_line_buffer[334]<=8'B11000000;oled_show_line_buffer[335]<=8'B01100000;oled_show_line_buffer[336]<=8'B00100000;oled_show_line_buffer[337]<=8'B00110000;oled_show_line_buffer[338]<=8'B00011000;oled_show_line_buffer[339]<=8'B00001100;oled_show_line_buffer[340]<=8'B00000100;end
                            10:begin oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[578]<=8'B00000001;oled_show_line_buffer[450]<=8'B10000000;oled_show_line_buffer[451]<=8'B10000000;oled_show_line_buffer[452]<=8'B11000000;oled_show_line_buffer[453]<=8'B01000000;oled_show_line_buffer[454]<=8'B01100000;oled_show_line_buffer[455]<=8'B00110000;oled_show_line_buffer[456]<=8'B00010000;oled_show_line_buffer[457]<=8'B00011000;oled_show_line_buffer[458]<=8'B00001000;oled_show_line_buffer[459]<=8'B00001100;oled_show_line_buffer[460]<=8'B00000110;oled_show_line_buffer[461]<=8'B00000010;oled_show_line_buffer[462]<=8'B00000011;oled_show_line_buffer[463]<=8'B00000001;oled_show_line_buffer[464]<=8'B00000001;oled_show_line_buffer[336]<=8'B10000000;oled_show_line_buffer[337]<=8'B10000000;oled_show_line_buffer[338]<=8'B11000000;oled_show_line_buffer[339]<=8'B01100000;oled_show_line_buffer[340]<=8'B00100000;end
                            11:begin oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[578]<=8'B00000001;oled_show_line_buffer[579]<=8'B00000001;oled_show_line_buffer[451]<=8'B10000000;oled_show_line_buffer[452]<=8'B10000000;oled_show_line_buffer[453]<=8'B11000000;oled_show_line_buffer[454]<=8'B01000000;oled_show_line_buffer[455]<=8'B01100000;oled_show_line_buffer[456]<=8'B00100000;oled_show_line_buffer[457]<=8'B00100000;oled_show_line_buffer[458]<=8'B00110000;oled_show_line_buffer[459]<=8'B00010000;oled_show_line_buffer[460]<=8'B00011000;oled_show_line_buffer[461]<=8'B00001000;oled_show_line_buffer[462]<=8'B00001100;oled_show_line_buffer[463]<=8'B00000100;oled_show_line_buffer[464]<=8'B00000110;oled_show_line_buffer[465]<=8'B00000010;oled_show_line_buffer[466]<=8'B00000010;oled_show_line_buffer[467]<=8'B00000011;oled_show_line_buffer[468]<=8'B00000001;oled_show_line_buffer[469]<=8'B00000001;oled_show_line_buffer[341]<=8'B10000000;oled_show_line_buffer[342]<=8'B10100000;end
                            12:begin oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[578]<=8'B00000001;oled_show_line_buffer[579]<=8'B00000001;oled_show_line_buffer[580]<=8'B00000001;oled_show_line_buffer[452]<=8'B10000000;oled_show_line_buffer[453]<=8'B10000000;oled_show_line_buffer[454]<=8'B10000000;oled_show_line_buffer[455]<=8'B11000000;oled_show_line_buffer[456]<=8'B01000000;oled_show_line_buffer[457]<=8'B01000000;oled_show_line_buffer[458]<=8'B01100000;oled_show_line_buffer[459]<=8'B00100000;oled_show_line_buffer[460]<=8'B00100000;oled_show_line_buffer[461]<=8'B00110000;oled_show_line_buffer[462]<=8'B00010000;oled_show_line_buffer[463]<=8'B00010000;oled_show_line_buffer[464]<=8'B00011000;oled_show_line_buffer[465]<=8'B00001000;oled_show_line_buffer[466]<=8'B00001000;oled_show_line_buffer[467]<=8'B00001000;oled_show_line_buffer[468]<=8'B00001100;oled_show_line_buffer[469]<=8'B00000100;oled_show_line_buffer[470]<=8'B00000100;oled_show_line_buffer[471]<=8'B00000110;oled_show_line_buffer[472]<=8'B00000010;end
                            13:begin oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[578]<=8'B00000011;oled_show_line_buffer[579]<=8'B00000001;oled_show_line_buffer[580]<=8'B00000001;oled_show_line_buffer[581]<=8'B00000001;oled_show_line_buffer[582]<=8'B00000001;oled_show_line_buffer[583]<=8'B00000001;oled_show_line_buffer[455]<=8'B10000000;oled_show_line_buffer[456]<=8'B10000000;oled_show_line_buffer[457]<=8'B10000000;oled_show_line_buffer[458]<=8'B10000000;oled_show_line_buffer[459]<=8'B11000000;oled_show_line_buffer[460]<=8'B01000000;oled_show_line_buffer[461]<=8'B01000000;oled_show_line_buffer[462]<=8'B01000000;oled_show_line_buffer[463]<=8'B01000000;oled_show_line_buffer[464]<=8'B01100000;oled_show_line_buffer[465]<=8'B00100000;oled_show_line_buffer[466]<=8'B00100000;oled_show_line_buffer[467]<=8'B00100000;oled_show_line_buffer[468]<=8'B00100000;oled_show_line_buffer[469]<=8'B00110000;oled_show_line_buffer[470]<=8'B00010000;oled_show_line_buffer[471]<=8'B00010000;end
                            14:begin oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[578]<=8'B00000010;oled_show_line_buffer[579]<=8'B00000010;oled_show_line_buffer[580]<=8'B00000011;oled_show_line_buffer[581]<=8'B00000001;oled_show_line_buffer[582]<=8'B00000001;oled_show_line_buffer[583]<=8'B00000001;oled_show_line_buffer[584]<=8'B00000001;oled_show_line_buffer[585]<=8'B00000001;oled_show_line_buffer[586]<=8'B00000001;oled_show_line_buffer[587]<=8'B00000001;oled_show_line_buffer[588]<=8'B00000001;oled_show_line_buffer[589]<=8'B00000001;oled_show_line_buffer[590]<=8'B00000001;oled_show_line_buffer[462]<=8'B10000000;oled_show_line_buffer[463]<=8'B10000000;oled_show_line_buffer[464]<=8'B10000000;oled_show_line_buffer[465]<=8'B10000000;oled_show_line_buffer[466]<=8'B10000000;oled_show_line_buffer[467]<=8'B10000000;oled_show_line_buffer[468]<=8'B10000000;oled_show_line_buffer[469]<=8'B10000000;oled_show_line_buffer[470]<=8'B10000000;oled_show_line_buffer[471]<=8'B11000000;oled_show_line_buffer[472]<=8'B01000000;oled_show_line_buffer[473]<=8'B01000000;oled_show_line_buffer[474]<=8'B01000000;oled_show_line_buffer[475]<=8'B01000000;oled_show_line_buffer[476]<=8'B01000000;end
                            15:begin oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[578]<=8'B00000001;oled_show_line_buffer[579]<=8'B00000001;oled_show_line_buffer[580]<=8'B00000001;oled_show_line_buffer[581]<=8'B00000001;oled_show_line_buffer[582]<=8'B00000001;oled_show_line_buffer[583]<=8'B00000001;oled_show_line_buffer[584]<=8'B00000001;oled_show_line_buffer[585]<=8'B00000001;oled_show_line_buffer[586]<=8'B00000001;oled_show_line_buffer[587]<=8'B00000001;oled_show_line_buffer[588]<=8'B00000001;oled_show_line_buffer[589]<=8'B00000001;oled_show_line_buffer[590]<=8'B00000001;oled_show_line_buffer[591]<=8'B00000001;oled_show_line_buffer[592]<=8'B00000001;oled_show_line_buffer[593]<=8'B00000001;oled_show_line_buffer[594]<=8'B00000001;oled_show_line_buffer[595]<=8'B00000001;oled_show_line_buffer[596]<=8'B00000001;oled_show_line_buffer[597]<=8'B00000001;oled_show_line_buffer[598]<=8'B00000001;oled_show_line_buffer[599]<=8'B00000001;oled_show_line_buffer[600]<=8'B00000001;oled_show_line_buffer[601]<=8'B00000001;end
                            16:begin oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[578]<=8'B00000001;oled_show_line_buffer[579]<=8'B00000001;oled_show_line_buffer[580]<=8'B00000001;oled_show_line_buffer[581]<=8'B00000001;oled_show_line_buffer[582]<=8'B00000001;oled_show_line_buffer[583]<=8'B00000001;oled_show_line_buffer[584]<=8'B00000001;oled_show_line_buffer[585]<=8'B00000011;oled_show_line_buffer[586]<=8'B00000010;oled_show_line_buffer[587]<=8'B00000010;oled_show_line_buffer[588]<=8'B00000010;oled_show_line_buffer[589]<=8'B00000010;oled_show_line_buffer[590]<=8'B00000010;oled_show_line_buffer[591]<=8'B00000010;oled_show_line_buffer[592]<=8'B00000010;oled_show_line_buffer[593]<=8'B00000010;oled_show_line_buffer[594]<=8'B00000110;oled_show_line_buffer[595]<=8'B00000100;oled_show_line_buffer[596]<=8'B00000100;oled_show_line_buffer[597]<=8'B00000100;oled_show_line_buffer[598]<=8'B00000100;oled_show_line_buffer[599]<=8'B00000100;oled_show_line_buffer[600]<=8'B00000100;oled_show_line_buffer[601]<=8'B00000100;oled_show_line_buffer[602]<=8'B00000100;oled_show_line_buffer[603]<=8'B00000100;oled_show_line_buffer[604]<=8'B00000101;end
                            17:begin oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[578]<=8'B00000001;oled_show_line_buffer[579]<=8'B00000001;oled_show_line_buffer[580]<=8'B00000011;oled_show_line_buffer[581]<=8'B00000010;oled_show_line_buffer[582]<=8'B00000010;oled_show_line_buffer[583]<=8'B00000010;oled_show_line_buffer[584]<=8'B00000110;oled_show_line_buffer[585]<=8'B00000100;oled_show_line_buffer[586]<=8'B00000100;oled_show_line_buffer[587]<=8'B00000100;oled_show_line_buffer[588]<=8'B00000100;oled_show_line_buffer[589]<=8'B00001100;oled_show_line_buffer[590]<=8'B00001000;oled_show_line_buffer[591]<=8'B00001000;oled_show_line_buffer[592]<=8'B00001000;oled_show_line_buffer[593]<=8'B00001000;oled_show_line_buffer[594]<=8'B00011000;oled_show_line_buffer[595]<=8'B00010000;oled_show_line_buffer[596]<=8'B00010000;oled_show_line_buffer[597]<=8'B00010000;oled_show_line_buffer[598]<=8'B00010000;oled_show_line_buffer[599]<=8'B00110000;oled_show_line_buffer[600]<=8'B00100000;oled_show_line_buffer[601]<=8'B00100000;oled_show_line_buffer[602]<=8'B00100000;oled_show_line_buffer[603]<=8'B00100000;end
                            18:begin oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[578]<=8'B00000011;oled_show_line_buffer[579]<=8'B00000010;oled_show_line_buffer[580]<=8'B00000010;oled_show_line_buffer[581]<=8'B00000110;oled_show_line_buffer[582]<=8'B00000100;oled_show_line_buffer[583]<=8'B00000100;oled_show_line_buffer[584]<=8'B00001100;oled_show_line_buffer[585]<=8'B00001000;oled_show_line_buffer[586]<=8'B00001000;oled_show_line_buffer[587]<=8'B00011000;oled_show_line_buffer[588]<=8'B00010000;oled_show_line_buffer[589]<=8'B00010000;oled_show_line_buffer[590]<=8'B00110000;oled_show_line_buffer[591]<=8'B00100000;oled_show_line_buffer[592]<=8'B00100000;oled_show_line_buffer[593]<=8'B01100000;oled_show_line_buffer[594]<=8'B01000000;oled_show_line_buffer[595]<=8'B01000000;oled_show_line_buffer[596]<=8'B01000000;oled_show_line_buffer[597]<=8'B11000000;oled_show_line_buffer[598]<=8'B10000000;oled_show_line_buffer[599]<=8'B10000000;oled_show_line_buffer[600]<=8'B10000000;end
                            19:begin oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[578]<=8'B00000010;oled_show_line_buffer[579]<=8'B00000110;oled_show_line_buffer[580]<=8'B00000100;oled_show_line_buffer[581]<=8'B00000100;oled_show_line_buffer[582]<=8'B00001100;oled_show_line_buffer[583]<=8'B00001000;oled_show_line_buffer[584]<=8'B00011000;oled_show_line_buffer[585]<=8'B00010000;oled_show_line_buffer[586]<=8'B00110000;oled_show_line_buffer[587]<=8'B00100000;oled_show_line_buffer[588]<=8'B01100000;oled_show_line_buffer[589]<=8'B01000000;oled_show_line_buffer[590]<=8'B01000000;oled_show_line_buffer[591]<=8'B11000000;oled_show_line_buffer[592]<=8'B10000000;oled_show_line_buffer[593]<=8'B10000000;oled_show_line_buffer[721]<=8'B00000001;oled_show_line_buffer[722]<=8'B00000001;oled_show_line_buffer[723]<=8'B00000011;oled_show_line_buffer[724]<=8'B00000010;oled_show_line_buffer[725]<=8'B00001110;oled_show_line_buffer[726]<=8'B00010100;oled_show_line_buffer[727]<=8'B00010100;oled_show_line_buffer[728]<=8'B00100100;end
                            20:begin oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[578]<=8'B00000110;oled_show_line_buffer[579]<=8'B00000100;oled_show_line_buffer[580]<=8'B00001100;oled_show_line_buffer[581]<=8'B00001000;oled_show_line_buffer[582]<=8'B00011000;oled_show_line_buffer[583]<=8'B00010000;oled_show_line_buffer[584]<=8'B00110000;oled_show_line_buffer[585]<=8'B01100000;oled_show_line_buffer[586]<=8'B01000000;oled_show_line_buffer[587]<=8'B11000000;oled_show_line_buffer[588]<=8'B10000000;oled_show_line_buffer[589]<=8'B10000000;oled_show_line_buffer[717]<=8'B00000001;oled_show_line_buffer[718]<=8'B00000001;oled_show_line_buffer[719]<=8'B00000011;oled_show_line_buffer[720]<=8'B00000110;oled_show_line_buffer[721]<=8'B00000100;oled_show_line_buffer[722]<=8'B00001100;oled_show_line_buffer[723]<=8'B00001000;oled_show_line_buffer[724]<=8'B00011000;oled_show_line_buffer[725]<=8'B00011000;oled_show_line_buffer[726]<=8'B00010000;end
                            21:begin oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[578]<=8'B00000110;oled_show_line_buffer[579]<=8'B00001100;oled_show_line_buffer[580]<=8'B00001000;oled_show_line_buffer[581]<=8'B00011000;oled_show_line_buffer[582]<=8'B00110000;oled_show_line_buffer[583]<=8'B01100000;oled_show_line_buffer[584]<=8'B01000000;oled_show_line_buffer[585]<=8'B11000000;oled_show_line_buffer[586]<=8'B10000000;oled_show_line_buffer[714]<=8'B00000001;oled_show_line_buffer[715]<=8'B00000011;oled_show_line_buffer[716]<=8'B00000010;oled_show_line_buffer[717]<=8'B00000110;oled_show_line_buffer[718]<=8'B00001100;oled_show_line_buffer[719]<=8'B00001000;oled_show_line_buffer[720]<=8'B00011000;oled_show_line_buffer[721]<=8'B00110000;oled_show_line_buffer[722]<=8'B01100000;oled_show_line_buffer[723]<=8'B01000000;oled_show_line_buffer[724]<=8'B01000000;end
                            22:begin oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[577]<=8'B00000111;oled_show_line_buffer[578]<=8'B00001100;oled_show_line_buffer[579]<=8'B00011000;oled_show_line_buffer[580]<=8'B00010000;oled_show_line_buffer[581]<=8'B00110000;oled_show_line_buffer[582]<=8'B01100000;oled_show_line_buffer[583]<=8'B11000000;oled_show_line_buffer[584]<=8'B10000000;oled_show_line_buffer[712]<=8'B00000001;oled_show_line_buffer[713]<=8'B00000011;oled_show_line_buffer[714]<=8'B00000110;oled_show_line_buffer[715]<=8'B00001100;oled_show_line_buffer[716]<=8'B00011000;oled_show_line_buffer[717]<=8'B00110000;oled_show_line_buffer[718]<=8'B00100000;oled_show_line_buffer[719]<=8'B01100000;oled_show_line_buffer[720]<=8'B11000000;oled_show_line_buffer[721]<=8'B10000000;oled_show_line_buffer[849]<=8'B00000001;oled_show_line_buffer[850]<=8'B00000011;oled_show_line_buffer[851]<=8'B10000010;end
                            23:begin oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[577]<=8'B00000111;oled_show_line_buffer[578]<=8'B00001100;oled_show_line_buffer[579]<=8'B00011000;oled_show_line_buffer[580]<=8'B01110000;oled_show_line_buffer[581]<=8'B11000000;oled_show_line_buffer[582]<=8'B10000000;oled_show_line_buffer[710]<=8'B00000001;oled_show_line_buffer[711]<=8'B00000011;oled_show_line_buffer[712]<=8'B00000110;oled_show_line_buffer[713]<=8'B00001100;oled_show_line_buffer[714]<=8'B00011000;oled_show_line_buffer[715]<=8'B00110000;oled_show_line_buffer[716]<=8'B01100000;oled_show_line_buffer[717]<=8'B11000000;oled_show_line_buffer[845]<=8'B10000001;oled_show_line_buffer[846]<=8'B00000011;oled_show_line_buffer[847]<=8'B00000110;oled_show_line_buffer[848]<=8'B00000100;end
                            24:begin oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000111;oled_show_line_buffer[577]<=8'B00001111;oled_show_line_buffer[578]<=8'B00011000;oled_show_line_buffer[579]<=8'B01110000;oled_show_line_buffer[580]<=8'B11000000;oled_show_line_buffer[581]<=8'B10000000;oled_show_line_buffer[709]<=8'B00000001;oled_show_line_buffer[710]<=8'B00000111;oled_show_line_buffer[711]<=8'B00001100;oled_show_line_buffer[712]<=8'B00111000;oled_show_line_buffer[713]<=8'B01100000;oled_show_line_buffer[714]<=8'B11000000;oled_show_line_buffer[715]<=8'B10000000;oled_show_line_buffer[843]<=8'B00000011;oled_show_line_buffer[844]<=8'B01000110;oled_show_line_buffer[845]<=8'B10001100;oled_show_line_buffer[846]<=8'B00011000;end
                            25:begin oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000111;oled_show_line_buffer[577]<=8'B00011111;oled_show_line_buffer[578]<=8'B01110000;oled_show_line_buffer[579]<=8'B11000000;oled_show_line_buffer[580]<=8'B10000000;oled_show_line_buffer[708]<=8'B00000011;oled_show_line_buffer[709]<=8'B00001110;oled_show_line_buffer[710]<=8'B00011000;oled_show_line_buffer[711]<=8'B01110000;oled_show_line_buffer[712]<=8'B11000000;oled_show_line_buffer[840]<=8'B00000001;oled_show_line_buffer[841]<=8'B00000111;oled_show_line_buffer[842]<=8'B00001100;oled_show_line_buffer[843]<=8'B00011000;end
                            26:begin oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[576]<=8'B00001111;oled_show_line_buffer[577]<=8'B00111011;oled_show_line_buffer[578]<=8'B11100000;oled_show_line_buffer[579]<=8'B10000000;oled_show_line_buffer[707]<=8'B00000111;oled_show_line_buffer[708]<=8'B00011100;oled_show_line_buffer[709]<=8'B01110000;oled_show_line_buffer[710]<=8'B11000000;oled_show_line_buffer[838]<=8'B00000001;oled_show_line_buffer[839]<=8'B00001111;oled_show_line_buffer[840]<=8'B00111000;oled_show_line_buffer[841]<=8'B01100000;end
                            27:begin oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[576]<=8'B00011111;oled_show_line_buffer[577]<=8'B11110011;oled_show_line_buffer[578]<=8'B10000000;oled_show_line_buffer[706]<=8'B00000111;oled_show_line_buffer[707]<=8'B00111100;oled_show_line_buffer[708]<=8'B11100000;oled_show_line_buffer[836]<=8'B00000001;oled_show_line_buffer[837]<=8'B00011111;oled_show_line_buffer[838]<=8'B11110000;oled_show_line_buffer[839]<=8'B10000000;oled_show_line_buffer[967]<=8'B00100001;end
                            28:begin oled_show_line_buffer[575]<=8'B00000111;oled_show_line_buffer[576]<=8'B11111111;oled_show_line_buffer[577]<=8'B10000011;oled_show_line_buffer[705]<=8'B00001111;oled_show_line_buffer[706]<=8'B11111000;oled_show_line_buffer[834]<=8'B00000001;oled_show_line_buffer[835]<=8'B00111111;oled_show_line_buffer[836]<=8'B11100000;end
                            29:begin oled_show_line_buffer[575]<=8'B00011111;oled_show_line_buffer[576]<=8'B11110011;oled_show_line_buffer[704]<=8'B01111111;oled_show_line_buffer[705]<=8'B11000000;oled_show_line_buffer[833]<=8'B11111111;oled_show_line_buffer[834]<=8'B10000000;oled_show_line_buffer[962]<=8'B01011111;end
                            30:begin oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[576]<=8'B11111111;oled_show_line_buffer[704]<=8'B11111111;oled_show_line_buffer[832]<=8'B11111111;oled_show_line_buffer[960]<=8'B01000011;end
                            31:begin oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[576]<=8'B11111111;oled_show_line_buffer[704]<=8'B00000011;oled_show_line_buffer[703]<=8'B11111110;oled_show_line_buffer[831]<=8'B00000111;oled_show_line_buffer[830]<=8'B11111100;oled_show_line_buffer[958]<=8'B01011111;end
                            32:begin oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[576]<=8'B00011111;oled_show_line_buffer[575]<=8'B11110011;oled_show_line_buffer[703]<=8'B00000001;oled_show_line_buffer[702]<=8'B00111111;oled_show_line_buffer[701]<=8'B11100000;oled_show_line_buffer[829]<=8'B00000111;oled_show_line_buffer[828]<=8'B11111100;oled_show_line_buffer[827]<=8'B10000000;oled_show_line_buffer[955]<=8'B00101111;end
                            33:begin oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[576]<=8'B00000111;oled_show_line_buffer[575]<=8'B00111111;oled_show_line_buffer[574]<=8'B11100000;oled_show_line_buffer[702]<=8'B00000001;oled_show_line_buffer[701]<=8'B00001111;oled_show_line_buffer[700]<=8'B01111000;oled_show_line_buffer[699]<=8'B11000000;oled_show_line_buffer[827]<=8'B00000011;oled_show_line_buffer[826]<=8'B00111110;oled_show_line_buffer[825]<=8'B11100000;oled_show_line_buffer[953]<=8'B00100001;end
                            34:begin oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[575]<=8'B00001111;oled_show_line_buffer[574]<=8'B01111000;oled_show_line_buffer[573]<=8'B11000000;oled_show_line_buffer[701]<=8'B00000001;oled_show_line_buffer[700]<=8'B00000111;oled_show_line_buffer[699]<=8'B00011100;oled_show_line_buffer[698]<=8'B11110000;oled_show_line_buffer[697]<=8'B10000000;oled_show_line_buffer[825]<=8'B00000011;oled_show_line_buffer[824]<=8'B00001110;oled_show_line_buffer[823]<=8'B00111000;oled_show_line_buffer[822]<=8'B11100000;oled_show_line_buffer[950]<=8'B00010001;end
                            35:begin oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[575]<=8'B00000111;oled_show_line_buffer[574]<=8'B00011100;oled_show_line_buffer[573]<=8'B01110000;oled_show_line_buffer[572]<=8'B11000000;oled_show_line_buffer[700]<=8'B00000001;oled_show_line_buffer[699]<=8'B00000011;oled_show_line_buffer[698]<=8'B00001110;oled_show_line_buffer[697]<=8'B00111000;oled_show_line_buffer[696]<=8'B11100000;oled_show_line_buffer[695]<=8'B10000000;oled_show_line_buffer[823]<=8'B00000001;oled_show_line_buffer[822]<=8'B00000111;oled_show_line_buffer[821]<=8'B00111100;oled_show_line_buffer[820]<=8'B01110000;end
                            36:begin oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[575]<=8'B00000111;oled_show_line_buffer[574]<=8'B00001100;oled_show_line_buffer[573]<=8'B00111000;oled_show_line_buffer[572]<=8'B01100000;oled_show_line_buffer[571]<=8'B11000000;oled_show_line_buffer[570]<=8'B10000000;oled_show_line_buffer[698]<=8'B00000011;oled_show_line_buffer[697]<=8'B00000110;oled_show_line_buffer[696]<=8'B00001100;oled_show_line_buffer[695]<=8'B00111000;oled_show_line_buffer[694]<=8'B01100000;oled_show_line_buffer[693]<=8'B11000000;oled_show_line_buffer[821]<=8'B00100001;oled_show_line_buffer[820]<=8'B01000011;oled_show_line_buffer[819]<=8'B10000110;oled_show_line_buffer[818]<=8'B10011100;end
                            37:begin oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[574]<=8'B00000110;oled_show_line_buffer[573]<=8'B00001100;oled_show_line_buffer[572]<=8'B00111000;oled_show_line_buffer[571]<=8'B01100000;oled_show_line_buffer[570]<=8'B11000000;oled_show_line_buffer[569]<=8'B10000000;oled_show_line_buffer[697]<=8'B00000001;oled_show_line_buffer[696]<=8'B00000011;oled_show_line_buffer[695]<=8'B00000110;oled_show_line_buffer[694]<=8'B00001100;oled_show_line_buffer[693]<=8'B00011000;oled_show_line_buffer[692]<=8'B00110000;oled_show_line_buffer[691]<=8'B11100000;oled_show_line_buffer[690]<=8'B10000000;oled_show_line_buffer[818]<=8'B10000001;oled_show_line_buffer[817]<=8'B00000011;oled_show_line_buffer[816]<=8'B00000110;oled_show_line_buffer[815]<=8'B00001100;end
                            38:begin oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[574]<=8'B00000110;oled_show_line_buffer[573]<=8'B00001100;oled_show_line_buffer[572]<=8'B00011000;oled_show_line_buffer[571]<=8'B00010000;oled_show_line_buffer[570]<=8'B00110000;oled_show_line_buffer[569]<=8'B01100000;oled_show_line_buffer[568]<=8'B11000000;oled_show_line_buffer[567]<=8'B10000000;oled_show_line_buffer[695]<=8'B00000001;oled_show_line_buffer[694]<=8'B00000011;oled_show_line_buffer[693]<=8'B00000110;oled_show_line_buffer[692]<=8'B00001100;oled_show_line_buffer[691]<=8'B00011000;oled_show_line_buffer[690]<=8'B00110000;oled_show_line_buffer[689]<=8'B00100000;oled_show_line_buffer[688]<=8'B01100000;oled_show_line_buffer[687]<=8'B11000000;oled_show_line_buffer[686]<=8'B10000000;oled_show_line_buffer[814]<=8'B10000001;end
                            39:begin oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[574]<=8'B00000011;oled_show_line_buffer[573]<=8'B00000110;oled_show_line_buffer[572]<=8'B00001100;oled_show_line_buffer[571]<=8'B00001000;oled_show_line_buffer[570]<=8'B00011000;oled_show_line_buffer[569]<=8'B00110000;oled_show_line_buffer[568]<=8'B01100000;oled_show_line_buffer[567]<=8'B01000000;oled_show_line_buffer[566]<=8'B11000000;oled_show_line_buffer[565]<=8'B10000000;oled_show_line_buffer[693]<=8'B00000001;oled_show_line_buffer[692]<=8'B00000001;oled_show_line_buffer[691]<=8'B00000011;oled_show_line_buffer[690]<=8'B00000110;oled_show_line_buffer[689]<=8'B00001100;oled_show_line_buffer[688]<=8'B00001000;oled_show_line_buffer[687]<=8'B00011000;oled_show_line_buffer[686]<=8'B00110000;oled_show_line_buffer[685]<=8'B01100000;oled_show_line_buffer[684]<=8'B01000000;end
                            40:begin oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[574]<=8'B00000011;oled_show_line_buffer[573]<=8'B00000010;oled_show_line_buffer[572]<=8'B00000110;oled_show_line_buffer[571]<=8'B00000100;oled_show_line_buffer[570]<=8'B00001100;oled_show_line_buffer[569]<=8'B00011000;oled_show_line_buffer[568]<=8'B00010000;oled_show_line_buffer[567]<=8'B00110000;oled_show_line_buffer[566]<=8'B00100000;oled_show_line_buffer[565]<=8'B01100000;oled_show_line_buffer[564]<=8'B11000000;oled_show_line_buffer[563]<=8'B10000000;oled_show_line_buffer[562]<=8'B10000000;oled_show_line_buffer[690]<=8'B00000001;oled_show_line_buffer[689]<=8'B00000001;oled_show_line_buffer[688]<=8'B00000011;oled_show_line_buffer[687]<=8'B00000010;oled_show_line_buffer[686]<=8'B00000110;oled_show_line_buffer[685]<=8'B00001100;oled_show_line_buffer[684]<=8'B00001000;end
                            41:begin oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[447]<=8'B10000000;oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[574]<=8'B00000001;oled_show_line_buffer[573]<=8'B00000011;oled_show_line_buffer[572]<=8'B00000010;oled_show_line_buffer[571]<=8'B00000110;oled_show_line_buffer[570]<=8'B00000100;oled_show_line_buffer[569]<=8'B00001100;oled_show_line_buffer[568]<=8'B00001000;oled_show_line_buffer[567]<=8'B00001000;oled_show_line_buffer[566]<=8'B00011000;oled_show_line_buffer[565]<=8'B00010000;oled_show_line_buffer[564]<=8'B00110000;oled_show_line_buffer[563]<=8'B00100000;oled_show_line_buffer[562]<=8'B01100000;oled_show_line_buffer[561]<=8'B01000000;oled_show_line_buffer[560]<=8'B11000000;oled_show_line_buffer[559]<=8'B10000000;oled_show_line_buffer[558]<=8'B10000000;oled_show_line_buffer[557]<=8'B10000000;oled_show_line_buffer[685]<=8'B00000001;oled_show_line_buffer[684]<=8'B00000001;oled_show_line_buffer[683]<=8'B00001011;oled_show_line_buffer[682]<=8'B00010010;end
                            42:begin oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[447]<=8'B10000000;oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[574]<=8'B00000001;oled_show_line_buffer[573]<=8'B00000001;oled_show_line_buffer[572]<=8'B00000011;oled_show_line_buffer[571]<=8'B00000010;oled_show_line_buffer[570]<=8'B00000010;oled_show_line_buffer[569]<=8'B00000110;oled_show_line_buffer[568]<=8'B00000100;oled_show_line_buffer[567]<=8'B00000100;oled_show_line_buffer[566]<=8'B00001100;oled_show_line_buffer[565]<=8'B00001000;oled_show_line_buffer[564]<=8'B00001000;oled_show_line_buffer[563]<=8'B00011000;oled_show_line_buffer[562]<=8'B00010000;oled_show_line_buffer[561]<=8'B00010000;oled_show_line_buffer[560]<=8'B00110000;oled_show_line_buffer[559]<=8'B00100000;oled_show_line_buffer[558]<=8'B00100000;oled_show_line_buffer[557]<=8'B00100000;oled_show_line_buffer[556]<=8'B01100000;oled_show_line_buffer[555]<=8'B01000000;oled_show_line_buffer[554]<=8'B01000000;oled_show_line_buffer[553]<=8'B11000000;oled_show_line_buffer[552]<=8'B10000000;end
                            43:begin oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[447]<=8'B10000000;oled_show_line_buffer[446]<=8'B10000000;oled_show_line_buffer[574]<=8'B00000001;oled_show_line_buffer[573]<=8'B00000001;oled_show_line_buffer[572]<=8'B00000001;oled_show_line_buffer[571]<=8'B00000001;oled_show_line_buffer[570]<=8'B00000001;oled_show_line_buffer[569]<=8'B00000011;oled_show_line_buffer[568]<=8'B00000010;oled_show_line_buffer[567]<=8'B00000010;oled_show_line_buffer[566]<=8'B00000010;oled_show_line_buffer[565]<=8'B00000110;oled_show_line_buffer[564]<=8'B00000100;oled_show_line_buffer[563]<=8'B00000100;oled_show_line_buffer[562]<=8'B00000100;oled_show_line_buffer[561]<=8'B00000100;oled_show_line_buffer[560]<=8'B00001100;oled_show_line_buffer[559]<=8'B00001000;oled_show_line_buffer[558]<=8'B00001000;oled_show_line_buffer[557]<=8'B00001000;oled_show_line_buffer[556]<=8'B00001000;oled_show_line_buffer[555]<=8'B00011000;oled_show_line_buffer[554]<=8'B00010000;oled_show_line_buffer[553]<=8'B00010000;end
                            44:begin oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[447]<=8'B10000000;oled_show_line_buffer[446]<=8'B10000000;oled_show_line_buffer[445]<=8'B10000000;oled_show_line_buffer[444]<=8'B10000000;oled_show_line_buffer[572]<=8'B00000001;oled_show_line_buffer[571]<=8'B00000001;oled_show_line_buffer[570]<=8'B00000001;oled_show_line_buffer[569]<=8'B00000001;oled_show_line_buffer[568]<=8'B00000001;oled_show_line_buffer[567]<=8'B00000001;oled_show_line_buffer[566]<=8'B00000001;oled_show_line_buffer[565]<=8'B00000001;oled_show_line_buffer[564]<=8'B00000001;oled_show_line_buffer[563]<=8'B00000001;oled_show_line_buffer[562]<=8'B00000011;oled_show_line_buffer[561]<=8'B00000010;oled_show_line_buffer[560]<=8'B00000010;oled_show_line_buffer[559]<=8'B00000010;oled_show_line_buffer[558]<=8'B00000010;oled_show_line_buffer[557]<=8'B00000010;oled_show_line_buffer[556]<=8'B00000010;oled_show_line_buffer[555]<=8'B00000010;oled_show_line_buffer[554]<=8'B00000010;oled_show_line_buffer[553]<=8'B00000110;oled_show_line_buffer[552]<=8'B00000100;oled_show_line_buffer[551]<=8'B00000100;oled_show_line_buffer[550]<=8'B00000101;oled_show_line_buffer[549]<=8'B00000101;oled_show_line_buffer[548]<=8'B00000101;end
                            45:begin oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[574]<=8'B00000001;oled_show_line_buffer[573]<=8'B00000001;oled_show_line_buffer[572]<=8'B00000001;oled_show_line_buffer[571]<=8'B00000001;oled_show_line_buffer[570]<=8'B00000001;oled_show_line_buffer[569]<=8'B00000001;oled_show_line_buffer[568]<=8'B00000001;oled_show_line_buffer[567]<=8'B00000001;oled_show_line_buffer[566]<=8'B00000001;oled_show_line_buffer[565]<=8'B00000001;oled_show_line_buffer[564]<=8'B00000001;oled_show_line_buffer[563]<=8'B00000001;oled_show_line_buffer[562]<=8'B00000001;oled_show_line_buffer[561]<=8'B00000001;oled_show_line_buffer[560]<=8'B00000001;oled_show_line_buffer[559]<=8'B00000001;oled_show_line_buffer[558]<=8'B00000001;oled_show_line_buffer[557]<=8'B00000001;oled_show_line_buffer[556]<=8'B00000001;oled_show_line_buffer[555]<=8'B00000001;oled_show_line_buffer[554]<=8'B00000001;oled_show_line_buffer[553]<=8'B00000001;oled_show_line_buffer[552]<=8'B00000001;oled_show_line_buffer[551]<=8'B00000001;end
                            46:begin oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[574]<=8'B00000001;oled_show_line_buffer[573]<=8'B00000001;oled_show_line_buffer[572]<=8'B00000001;oled_show_line_buffer[571]<=8'B00000001;oled_show_line_buffer[570]<=8'B00000001;oled_show_line_buffer[569]<=8'B00000001;oled_show_line_buffer[568]<=8'B00000001;oled_show_line_buffer[567]<=8'B00000001;oled_show_line_buffer[439]<=8'B10000000;oled_show_line_buffer[438]<=8'B10000000;oled_show_line_buffer[437]<=8'B10000000;oled_show_line_buffer[436]<=8'B10000000;oled_show_line_buffer[435]<=8'B10000000;oled_show_line_buffer[434]<=8'B10000000;oled_show_line_buffer[433]<=8'B10000000;oled_show_line_buffer[432]<=8'B10000000;oled_show_line_buffer[431]<=8'B10000000;oled_show_line_buffer[430]<=8'B11000000;oled_show_line_buffer[429]<=8'B01000000;oled_show_line_buffer[428]<=8'B01000000;oled_show_line_buffer[427]<=8'B01000000;oled_show_line_buffer[426]<=8'B01000000;oled_show_line_buffer[425]<=8'B01000000;oled_show_line_buffer[424]<=8'B01000000;oled_show_line_buffer[423]<=8'B01000000;oled_show_line_buffer[422]<=8'B01000000;oled_show_line_buffer[421]<=8'B01000000;oled_show_line_buffer[420]<=8'B01000000;end
                            47:begin oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[574]<=8'B00000001;oled_show_line_buffer[573]<=8'B00000001;oled_show_line_buffer[572]<=8'B00000001;oled_show_line_buffer[444]<=8'B10000000;oled_show_line_buffer[443]<=8'B10000000;oled_show_line_buffer[442]<=8'B10000000;oled_show_line_buffer[441]<=8'B10000000;oled_show_line_buffer[440]<=8'B11000000;oled_show_line_buffer[439]<=8'B01000000;oled_show_line_buffer[438]<=8'B01000000;oled_show_line_buffer[437]<=8'B01000000;oled_show_line_buffer[436]<=8'B01000000;oled_show_line_buffer[435]<=8'B01100000;oled_show_line_buffer[434]<=8'B00100000;oled_show_line_buffer[433]<=8'B00100000;oled_show_line_buffer[432]<=8'B00100000;oled_show_line_buffer[431]<=8'B00100000;oled_show_line_buffer[430]<=8'B00110000;oled_show_line_buffer[429]<=8'B00010000;oled_show_line_buffer[428]<=8'B00010000;oled_show_line_buffer[427]<=8'B00010000;oled_show_line_buffer[426]<=8'B00010000;oled_show_line_buffer[425]<=8'B00011000;oled_show_line_buffer[424]<=8'B00001000;oled_show_line_buffer[423]<=8'B00001000;oled_show_line_buffer[422]<=8'B00001000;oled_show_line_buffer[421]<=8'B00001000;end
                            48:begin oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[574]<=8'B00000001;oled_show_line_buffer[446]<=8'B10000000;oled_show_line_buffer[445]<=8'B10000000;oled_show_line_buffer[444]<=8'B10000000;oled_show_line_buffer[443]<=8'B11000000;oled_show_line_buffer[442]<=8'B01000000;oled_show_line_buffer[441]<=8'B01000000;oled_show_line_buffer[440]<=8'B01100000;oled_show_line_buffer[439]<=8'B00100000;oled_show_line_buffer[438]<=8'B00100000;oled_show_line_buffer[437]<=8'B00110000;oled_show_line_buffer[436]<=8'B00010000;oled_show_line_buffer[435]<=8'B00010000;oled_show_line_buffer[434]<=8'B00011000;oled_show_line_buffer[433]<=8'B00001000;oled_show_line_buffer[432]<=8'B00001000;oled_show_line_buffer[431]<=8'B00001100;oled_show_line_buffer[430]<=8'B00000100;oled_show_line_buffer[429]<=8'B00000100;oled_show_line_buffer[428]<=8'B00000100;oled_show_line_buffer[427]<=8'B00000110;oled_show_line_buffer[426]<=8'B00000010;oled_show_line_buffer[425]<=8'B00000010;oled_show_line_buffer[424]<=8'B00000010;end
                            49:begin oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[447]<=8'B10000000;oled_show_line_buffer[446]<=8'B10000000;oled_show_line_buffer[445]<=8'B11000000;oled_show_line_buffer[444]<=8'B01000000;oled_show_line_buffer[443]<=8'B01000000;oled_show_line_buffer[442]<=8'B01100000;oled_show_line_buffer[441]<=8'B00100000;oled_show_line_buffer[440]<=8'B00110000;oled_show_line_buffer[439]<=8'B00010000;oled_show_line_buffer[438]<=8'B00011000;oled_show_line_buffer[437]<=8'B00001000;oled_show_line_buffer[436]<=8'B00001100;oled_show_line_buffer[435]<=8'B00000100;oled_show_line_buffer[434]<=8'B00000100;oled_show_line_buffer[433]<=8'B00000110;oled_show_line_buffer[432]<=8'B00000010;oled_show_line_buffer[431]<=8'B00000011;oled_show_line_buffer[430]<=8'B00000001;oled_show_line_buffer[429]<=8'B00000001;oled_show_line_buffer[301]<=8'B10000000;oled_show_line_buffer[300]<=8'B10000000;oled_show_line_buffer[299]<=8'B11010000;oled_show_line_buffer[298]<=8'B01001000;oled_show_line_buffer[297]<=8'B01001000;oled_show_line_buffer[296]<=8'B01000100;end
                            50:begin oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[575]<=8'B00000011;oled_show_line_buffer[447]<=8'B10000000;oled_show_line_buffer[446]<=8'B11000000;oled_show_line_buffer[445]<=8'B01000000;oled_show_line_buffer[444]<=8'B01100000;oled_show_line_buffer[443]<=8'B00100000;oled_show_line_buffer[442]<=8'B00110000;oled_show_line_buffer[441]<=8'B00010000;oled_show_line_buffer[440]<=8'B00011000;oled_show_line_buffer[439]<=8'B00001100;oled_show_line_buffer[438]<=8'B00000100;oled_show_line_buffer[437]<=8'B00000110;oled_show_line_buffer[436]<=8'B00000010;oled_show_line_buffer[435]<=8'B00000011;oled_show_line_buffer[434]<=8'B00000001;oled_show_line_buffer[433]<=8'B00000001;oled_show_line_buffer[305]<=8'B10000000;oled_show_line_buffer[304]<=8'B11000000;oled_show_line_buffer[303]<=8'B01000000;oled_show_line_buffer[302]<=8'B01100000;oled_show_line_buffer[301]<=8'B00100000;oled_show_line_buffer[300]<=8'B00110000;oled_show_line_buffer[299]<=8'B00010000;oled_show_line_buffer[298]<=8'B00011000;end
                            51:begin oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[447]<=8'B10000000;oled_show_line_buffer[446]<=8'B11000000;oled_show_line_buffer[445]<=8'B01100000;oled_show_line_buffer[444]<=8'B00100000;oled_show_line_buffer[443]<=8'B00110000;oled_show_line_buffer[442]<=8'B00011000;oled_show_line_buffer[441]<=8'B00001100;oled_show_line_buffer[440]<=8'B00000100;oled_show_line_buffer[439]<=8'B00000110;oled_show_line_buffer[438]<=8'B00000011;oled_show_line_buffer[437]<=8'B00000001;oled_show_line_buffer[309]<=8'B10000000;oled_show_line_buffer[308]<=8'B10000000;oled_show_line_buffer[307]<=8'B11000000;oled_show_line_buffer[306]<=8'B01100000;oled_show_line_buffer[305]<=8'B00100000;oled_show_line_buffer[304]<=8'B00110000;oled_show_line_buffer[303]<=8'B00011000;oled_show_line_buffer[302]<=8'B00001100;oled_show_line_buffer[301]<=8'B00000100;oled_show_line_buffer[300]<=8'B00000100;end
                            52:begin oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[447]<=8'B11000000;oled_show_line_buffer[446]<=8'B01100000;oled_show_line_buffer[445]<=8'B00110000;oled_show_line_buffer[444]<=8'B00010000;oled_show_line_buffer[443]<=8'B00011000;oled_show_line_buffer[442]<=8'B00001100;oled_show_line_buffer[441]<=8'B00000110;oled_show_line_buffer[440]<=8'B00000011;oled_show_line_buffer[439]<=8'B00000001;oled_show_line_buffer[311]<=8'B10000000;oled_show_line_buffer[310]<=8'B11000000;oled_show_line_buffer[309]<=8'B01100000;oled_show_line_buffer[308]<=8'B00110000;oled_show_line_buffer[307]<=8'B00011000;oled_show_line_buffer[306]<=8'B00001000;oled_show_line_buffer[305]<=8'B00001100;oled_show_line_buffer[304]<=8'B00000110;oled_show_line_buffer[303]<=8'B00000011;oled_show_line_buffer[302]<=8'B00000001;oled_show_line_buffer[174]<=8'B10000001;oled_show_line_buffer[173]<=8'B10000001;end
                            53:begin oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[448]<=8'B10000000;oled_show_line_buffer[447]<=8'B11000000;oled_show_line_buffer[446]<=8'B01100000;oled_show_line_buffer[445]<=8'B00110000;oled_show_line_buffer[444]<=8'B00011100;oled_show_line_buffer[443]<=8'B00000110;oled_show_line_buffer[442]<=8'B00000011;oled_show_line_buffer[441]<=8'B00000001;oled_show_line_buffer[313]<=8'B10000000;oled_show_line_buffer[312]<=8'B11000000;oled_show_line_buffer[311]<=8'B01100000;oled_show_line_buffer[310]<=8'B00110000;oled_show_line_buffer[309]<=8'B00011000;oled_show_line_buffer[308]<=8'B00001100;oled_show_line_buffer[307]<=8'B00000111;oled_show_line_buffer[306]<=8'B00000001;oled_show_line_buffer[178]<=8'B10000000;oled_show_line_buffer[177]<=8'B11000000;oled_show_line_buffer[176]<=8'B01000000;end
                            54:begin oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[448]<=8'B11000000;oled_show_line_buffer[447]<=8'B11100000;oled_show_line_buffer[446]<=8'B00110000;oled_show_line_buffer[445]<=8'B00011100;oled_show_line_buffer[444]<=8'B00000110;oled_show_line_buffer[443]<=8'B00000011;oled_show_line_buffer[442]<=8'B00000001;oled_show_line_buffer[314]<=8'B11000000;oled_show_line_buffer[313]<=8'B01100000;oled_show_line_buffer[312]<=8'B00111000;oled_show_line_buffer[311]<=8'B00001100;oled_show_line_buffer[310]<=8'B00000110;oled_show_line_buffer[309]<=8'B00000011;oled_show_line_buffer[181]<=8'B10000100;oled_show_line_buffer[180]<=8'B11000011;oled_show_line_buffer[179]<=8'B01100000;oled_show_line_buffer[178]<=8'B00110000;end
                            55:begin oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[576]<=8'B00000011;oled_show_line_buffer[448]<=8'B11000000;oled_show_line_buffer[447]<=8'B11110000;oled_show_line_buffer[446]<=8'B00011100;oled_show_line_buffer[445]<=8'B00000110;oled_show_line_buffer[444]<=8'B00000011;oled_show_line_buffer[316]<=8'B10000000;oled_show_line_buffer[315]<=8'B11100000;oled_show_line_buffer[314]<=8'B00110000;oled_show_line_buffer[313]<=8'B00011100;oled_show_line_buffer[312]<=8'B00000111;oled_show_line_buffer[311]<=8'B00000001;oled_show_line_buffer[183]<=8'B11000000;oled_show_line_buffer[182]<=8'B01100000;oled_show_line_buffer[181]<=8'B00110100;end
                            56:begin oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[449]<=8'B10000000;oled_show_line_buffer[448]<=8'B11100000;oled_show_line_buffer[447]<=8'B10111000;oled_show_line_buffer[446]<=8'B00001110;oled_show_line_buffer[445]<=8'B00000011;oled_show_line_buffer[317]<=8'B11000000;oled_show_line_buffer[316]<=8'B01110000;oled_show_line_buffer[315]<=8'B00011100;oled_show_line_buffer[314]<=8'B00000111;oled_show_line_buffer[313]<=8'B00000001;oled_show_line_buffer[185]<=8'B11100000;oled_show_line_buffer[184]<=8'B00111000;oled_show_line_buffer[183]<=8'B00001100;end
                            57:begin oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[449]<=8'B10000000;oled_show_line_buffer[448]<=8'B11110000;oled_show_line_buffer[447]<=8'B10011110;oled_show_line_buffer[446]<=8'B00000011;oled_show_line_buffer[318]<=8'B11000000;oled_show_line_buffer[317]<=8'B01111000;oled_show_line_buffer[316]<=8'B00001111;oled_show_line_buffer[315]<=8'B00000001;oled_show_line_buffer[187]<=8'B11110000;oled_show_line_buffer[186]<=8'B00011110;oled_show_line_buffer[185]<=8'B00000011;end
                            58:begin oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[449]<=8'B11000000;oled_show_line_buffer[448]<=8'B11111110;oled_show_line_buffer[447]<=8'B10000011;oled_show_line_buffer[319]<=8'B11100000;oled_show_line_buffer[318]<=8'B00111111;oled_show_line_buffer[317]<=8'B00000001;oled_show_line_buffer[189]<=8'B11111000;oled_show_line_buffer[188]<=8'B00001110;end
                            59:begin oled_show_line_buffer[577]<=8'B00000011;oled_show_line_buffer[449]<=8'B11110000;oled_show_line_buffer[448]<=8'B10011111;oled_show_line_buffer[320]<=8'B11111100;oled_show_line_buffer[319]<=8'B00000111;oled_show_line_buffer[191]<=8'B11111110;oled_show_line_buffer[190]<=8'B00000011;oled_show_line_buffer[62]<=8'B11110010;end
                            endcase
                            
                            //oled_show_line_buffer[574]<=8'B00000100;oled_show_line_buffer[573]<=8'B00001000;oled_show_line_buffer[572]<=8'B00001000;oled_show_line_buffer[571]<=8'B00010000;oled_show_line_buffer[570]<=8'B00100000;oled_show_line_buffer[569]<=8'B00100000;oled_show_line_buffer[568]<=8'B01000000;oled_show_line_buffer[567]<=8'B10000000;oled_show_line_buffer[694]<=8'B00000001;oled_show_line_buffer[693]<=8'B00000001;oled_show_line_buffer[692]<=8'B00000010;oled_show_line_buffer[691]<=8'B00000100;oled_show_line_buffer[690]<=8'B00001000;oled_show_line_buffer[689]<=8'B00001000;oled_show_line_buffer[688]<=8'B00010000;oled_show_line_buffer[687]<=8'B00100000;oled_show_line_buffer[686]<=8'B00100000;oled_show_line_buffer[685]<=8'B01000000;oled_show_line_buffer[684]<=8'B10000000;oled_show_line_buffer[811]<=8'B00000001;oled_show_line_buffer[810]<=8'B00000001;
                        end
                    endcase
                end
            DRAW:begin
                if(send_done)begin
                    if(draw_st==DRAW_INIT_FINISHED)
                            counter<=counter+1;
                    case(draw_st)
                        DRAW_INIT1:draw_st<=DRAW_INIT2;
                        DRAW_INIT2:draw_st<=DRAW_INIT3;
                        DRAW_INIT3:draw_st<=DRAW_INIT_FINISHED;
                        DRAW_INIT_FINISHED:begin
                            if(counter%128==0)draw_st<=DRAW_INIT1;
                        end
                    endcase
                end
                if(counter==8*128-1)begin
                    cur_st<=FINISH;
                end
            end
            FINISH:begin
                if(show_st==DRAW_CLOCK)begin
                    cur_st<=WAITE;
                    show_st<=DRAW_LINE;
                    for(i=0;i<1024;i=i+1)begin
                        oled_show_line_buffer[i]<=oled_show_buffer[i];
                    end
                end
                else if(show_st==DRAW_LINE)begin
                    cur_st<=WAITE;
                    show_st<=DRAW_CLOCK;
                end
            end
        endcase
    end

    always@(*)begin
        case(cur_st)
            WAITE:begin spi_send=0;spi_data=0; end
            DRAW:begin 
                spi_send=1;
                case(draw_st)
                    DRAW_INIT1:begin spi_data=8'hb0 | (counter/128);dc=0;end
                    DRAW_INIT2:begin spi_data=8'h10;dc=0;end
                    DRAW_INIT3:begin spi_data=8'h00;dc=0;end
                    DRAW_INIT_FINISHED:begin spi_data=oled_show_line_buffer[counter];dc=1;end
                    default:begin spi_data=0; end
                endcase
            end
            FINISH:begin spi_send=0;spi_data=0; end
            default:begin spi_send=0;spi_data=0; end
        endcase
    end

endmodule
