/**
 * @module bin2bcd
 * @brief Converts a binary number to binary-coded decimal (BCD) representation.
 *
 * This module takes a binary input and converts it to BCD format. The BCD output
 * consists of separate digits representing thousands, hundreds, tens, and ones.
 *
 * @param W The width of the input binary number.
 * @param bin The binary input to be converted to BCD.
 * @param bcd The BCD output representing the converted binary number.
 */
module bin2bcd #(
    parameter W = 18  // input width
) (
    input      [    W-1 : 0] bin,  // binary
    output reg [W+(W-4)/3:0] bcd   // bcd {...,thousands,hundreds,tens,ones}
);

  integer i, j;

  always @(bin) begin
    for (i = 0; i <= W + (W - 4) / 3; i = i + 1) bcd[i] = 0;  // initialize with zeros
    bcd[W-1:0] = bin;  // initialize with input vector
    for (i = 0; i <= W - 4; i = i + 1)  // iterate on structure depth
      for (j = 0; j <= i / 3; j = j + 1)  // iterate on structure width
        if (bcd[W-i+4*j-:4] > 4)  // if > 4
          bcd[W-i+4*j-:4] = bcd[W-i+4*j-:4] + 4'd3;  // add 3
  end

endmodule
