`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/08/25 09:40:00
// Design Name: 
// Module Name: unixCounter
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module unixCounter #(
    parameter N = 64,  //计数器位数
    parameter M = 26   //分频计数器位数
) (
    input wire clk,
    input wire reset_n,
    input wire load_n,
    input wire go,
    input wire [N-1:0] set_counter,
    output reg [N-1:0] counter
);
  reg [M-1:0] division_counter;
  wire clk1Hz;
  //localparam divisionM=50000000;
  localparam divisionM = 5;
  initial begin
    division_counter = 64'b0;
    counter = 64'b1;
  end


  //分频计数器加
  always @(posedge clk) begin
    if (!reset_n) begin
      counter <= 0;
      division_counter <= 0;
    end else if (!load_n) begin
      counter <= set_counter;
      division_counter <= 0;
    end else if (go)
      if (division_counter < divisionM) division_counter <= division_counter + 1;
      else division_counter <= 0;
  end


  assign clk1Hz = (division_counter == divisionM) ? 1'b1 : 1'b0;

  //1Hz上升沿
  always @(posedge clk1Hz) counter <= counter + 1;

endmodule
